LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY MBE IS
PORT (A_SIG, B_SIG : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      OUT_MULT : OUT STD_LOGIC_VECTOR (63 DOWNTO 0));
END ENTITY;

ARCHITECTURE beh OF MBE IS

COMPONENT HA IS
PORT (input1, input2 : IN STD_LOGIC;
      out_HA : OUT STD_LOGIC;
      carry_out : OUT STD_LOGIC);
END COMPONENT;

COMPONENT FA IS
PORT (input1, input2 : IN STD_LOGIC;
      carry_in : IN STD_LOGIC;
      out_FA : OUT STD_LOGIC;
      carry_out : OUT STD_LOGIC);
END COMPONENT;

COMPONENT MUX_PRODUCT IS
PORT (IN1, IN2, IN3 : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
      SELECTOR : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      OUT_MUX : OUT STD_LOGIC_VECTOR (32 DOWNTO 0));
END COMPONENT;

SIGNAL A2, A, ZEROS : STD_LOGIC_VECTOR (32 DOWNTO 0);

SIGNAL SELECTOR_TABLE_0, SELECTOR_TABLE_1, SELECTOR_TABLE_2, SELECTOR_TABLE_3, SELECTOR_TABLE_4
     , SELECTOR_TABLE_5, SELECTOR_TABLE_6, SELECTOR_TABLE_7, SELECTOR_TABLE_8, SELECTOR_TABLE_9
     , SELECTOR_TABLE_10, SELECTOR_TABLE_11, SELECTOR_TABLE_12, SELECTOR_TABLE_13, SELECTOR_TABLE_14, 
       SELECTOR_TABLE_15, SELECTOR_TABLE_16 : STD_LOGIC_VECTOR (2 DOWNTO 0);

SIGNAL OUT_MUX_0, OUT_MUX_1, OUT_MUX_2, OUT_MUX_3, OUT_MUX_4, OUT_MUX_5, OUT_MUX_6, OUT_MUX_7, OUT_MUX_8,
       OUT_MUX_9, OUT_MUX_10, OUT_MUX_11, OUT_MUX_12, OUT_MUX_13, OUT_MUX_14, OUT_MUX_15, OUT_MUX_16 : STD_LOGIC_VECTOR (32 DOWNTO 0);

--PARTIAL PRODUCT INITIAL STRUCTURE
SIGNAL PP0, PP1, PP2,PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, 
       PP11, PP12, PP13, PP14, PP15, PP16 : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0'); 

--PARTIAL PRODUCT 1th LEVEL (TRIANGLE STRUCTURE)
SIGNAL PARTIAL_PRODUCT_0, PARTIAL_PRODUCT_1, PARTIAL_PRODUCT_2,PARTIAL_PRODUCT_3, PARTIAL_PRODUCT_4, 
       PARTIAL_PRODUCT_5, PARTIAL_PRODUCT_6, PARTIAL_PRODUCT_7, PARTIAL_PRODUCT_8, PARTIAL_PRODUCT_9, PARTIAL_PRODUCT_10, 
       PARTIAL_PRODUCT_11, PARTIAL_PRODUCT_12, PARTIAL_PRODUCT_13, PARTIAL_PRODUCT_14, PARTIAL_PRODUCT_15, PARTIAL_PRODUCT_16 : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0');

--PARTIAL PRODUCT 2th LEVEL --> PARTIAL_PRODUCT_i_1
SIGNAL PARTIAL_PRODUCT_0_1, PARTIAL_PRODUCT_1_1, PARTIAL_PRODUCT_2_1,PARTIAL_PRODUCT_3_1, 
       PARTIAL_PRODUCT_4_1, PARTIAL_PRODUCT_5_1, PARTIAL_PRODUCT_6_1, PARTIAL_PRODUCT_7_1, 
       PARTIAL_PRODUCT_8_1, PARTIAL_PRODUCT_9_1, PARTIAL_PRODUCT_10_1, PARTIAL_PRODUCT_11_1,
       PARTIAL_PRODUCT_12_1 : STD_LOGIC_VECTOR (63 DOWNTO 0) := (OTHERS =>'0');
  

--PARTIAL PRODUCT 3th LEVEL --> PARTIAL_PRODUCT_i_2
SIGNAL PARTIAL_PRODUCT_0_2,PARTIAL_PRODUCT_1_2,PARTIAL_PRODUCT_2_2, PARTIAL_PRODUCT_3_2, PARTIAL_PRODUCT_4_2,
       PARTIAL_PRODUCT_5_2, PARTIAL_PRODUCT_6_2, PARTIAL_PRODUCT_7_2, PARTIAL_PRODUCT_8_2 : STD_LOGIC_VECTOR (63 DOWNTO 0) := (OTHERS =>'0');

--PARTIAL PRODUCT 4th LEVEL --> PARTIAL_PRODUCT_i_3
SIGNAL PARTIAL_PRODUCT_0_3, PARTIAL_PRODUCT_1_3, PARTIAL_PRODUCT_2_3, PARTIAL_PRODUCT_3_3, PARTIAL_PRODUCT_4_3, PARTIAL_PRODUCT_5_3,
       PARTIAL_PRODUCT_6_3, PARTIAL_PRODUCT_7_3, PARTIAL_PRODUCT_8_3 : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0');

--PARTIAL PRODUCT 5th LEVEL --> PARTIAL_PRODUCT_i_4
SIGNAL PARTIAL_PRODUCT_0_4, PARTIAL_PRODUCT_1_4, PARTIAL_PRODUCT_2_4, PARTIAL_PRODUCT_3_4, PARTIAL_PRODUCT_4_4, PARTIAL_PRODUCT_5_4 : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0');

--PARTIAL PRODUCT 6th LEVEL --> PARTIAL_PRODUCT_i_5
SIGNAL PARTIAL_PRODUCT_0_5, PARTIAL_PRODUCT_1_5, PARTIAL_PRODUCT_2_5, PARTIAL_PRODUCT_3_5: STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0');

--PARTIAL PRODUCT 7TH LEVEL -->PARTIAL_PRODUCT_i_6
SIGNAL PARTIAL_PRODUCT_0_6, PARTIAL_PRODUCT_1_6,PARTIAL_PRODUCT_0_7, CARRY_OUT_7 : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS =>'0');
SIGNAL CARRY_6 :STD_LOGIC;

BEGIN

A(32) <= '0'; A(31 DOWNTO 0) <= A_SIG;
A2(32 DOWNTO 1) <= A_SIG; A2(0) <='0';
ZEROS <= (others => '0');



--DEFINE SELECTOR_TABLE_i
SELECTOR_TABLE_0 <= B_SIG(1 DOWNTO 0) & '0';
SELECTOR_TABLE_1 <= B_SIG(3 DOWNTO 1);
SELECTOR_TABLE_2 <= B_SIG(5 DOWNTO 3);
SELECTOR_TABLE_3 <= B_SIG(7 DOWNTO 5);
SELECTOR_TABLE_4 <= B_SIG(9 DOWNTO 7);
SELECTOR_TABLE_5 <= B_SIG(11 DOWNTO 9);
SELECTOR_TABLE_6 <= B_SIG(13 DOWNTO 11);
SELECTOR_TABLE_7 <= B_SIG(15 DOWNTO 13);
SELECTOR_TABLE_8 <= B_SIG(17 DOWNTO 15);
SELECTOR_TABLE_9 <= B_SIG(19 DOWNTO 17);
SELECTOR_TABLE_10 <= B_SIG(21 DOWNTO 19);
SELECTOR_TABLE_11 <= B_SIG(23 DOWNTO 21);
SELECTOR_TABLE_12 <= B_SIG(25 DOWNTO 23);
SELECTOR_TABLE_13 <= B_SIG(27 DOWNTO 25);
SELECTOR_TABLE_14 <= B_SIG(29 DOWNTO 27);
SELECTOR_TABLE_15 <= B_SIG(31 DOWNTO 29);
SELECTOR_TABLE_16 <= "00" & B_SIG(31);

--MUX SELECTOR POSITIVE PARTIAL PRODUCT
MUX_PRODUCT_0 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_0, OUT_MUX_0);
MUX_PRODUCT_1 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_1, OUT_MUX_1);
MUX_PRODUCT_2 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_2, OUT_MUX_2);
MUX_PRODUCT_3 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_3, OUT_MUX_3);
MUX_PRODUCT_4 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_4, OUT_MUX_4);
MUX_PRODUCT_5 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_5, OUT_MUX_5);
MUX_PRODUCT_6 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_6, OUT_MUX_6);
MUX_PRODUCT_7 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_7,OUT_MUX_7);
MUX_PRODUCT_8 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_8, OUT_MUX_8);
MUX_PRODUCT_9 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_9, OUT_MUX_9);
MUX_PRODUCT_10 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_10, OUT_MUX_10);
MUX_PRODUCT_11 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_11, OUT_MUX_11);
MUX_PRODUCT_12 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_12, OUT_MUX_12);
MUX_PRODUCT_13 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_13, OUT_MUX_13);
MUX_PRODUCT_14 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_14, OUT_MUX_14);
MUX_PRODUCT_15 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_15, OUT_MUX_15);
MUX_PRODUCT_16 : MUX_PRODUCT PORT MAP (ZEROS, A, A2,SELECTOR_TABLE_16, OUT_MUX_16);

--PARTIAL PRODUCT GENERATION (POSITIVE AND NEGATIVE)
PP0(32 DOWNTO 0)<= OUT_MUX_0 WHEN SELECTOR_TABLE_0(2)='0' ELSE NOT(OUT_MUX_0);
PP0 (34 DOWNTO 33) <= (OTHERS => SELECTOR_TABLE_0(2));
PP0 (35) <= NOT (SELECTOR_TABLE_0(2));

PP1(34 DOWNTO 2) <= OUT_MUX_1 WHEN SELECTOR_TABLE_1(2)='0' ELSE NOT(OUT_MUX_1);
PP1(0) <= SELECTOR_TABLE_0(2);
PP1(36) <= '1'; PP1(35) <= NOT (SELECTOR_TABLE_1(2));

PP2(36 DOWNTO 4) <= OUT_MUX_2 WHEN SELECTOR_TABLE_2(2)='0' ELSE NOT(OUT_MUX_2);
PP2(2) <= SELECTOR_TABLE_1(2);
PP2(38) <= '1'; PP2(37) <= NOT (SELECTOR_TABLE_2(2));

PP3(38 DOWNTO 6) <= OUT_MUX_3 WHEN SELECTOR_TABLE_3(2)='0' ELSE NOT(OUT_MUX_3);
PP3(4) <= SELECTOR_TABLE_2(2);
PP3(40) <= '1'; PP3(39) <= NOT (SELECTOR_TABLE_3(2));

PP4(40 DOWNTO 8) <= OUT_MUX_4 WHEN SELECTOR_TABLE_4(2)='0' ELSE NOT(OUT_MUX_4);
PP4(6) <= SELECTOR_TABLE_3(2); --PREC
PP4(42) <= '1'; PP4(41) <= NOT (SELECTOR_TABLE_4(2));

PP5(42 DOWNTO 10) <= OUT_MUX_5 WHEN SELECTOR_TABLE_5(2)='0' ELSE NOT(OUT_MUX_5);
PP5(8) <= SELECTOR_TABLE_4(2); --PREC
PP5(44) <= '1'; PP5(43) <= NOT (SELECTOR_TABLE_5(2));

PP6(44 DOWNTO 12) <= OUT_MUX_6 WHEN SELECTOR_TABLE_6(2)='0' ELSE NOT(OUT_MUX_6);
PP6(10) <= SELECTOR_TABLE_5(2); --PREC
PP6(46) <= '1'; PP6(45) <= NOT (SELECTOR_TABLE_6(2));

PP7(46 DOWNTO 14) <= OUT_MUX_7 WHEN SELECTOR_TABLE_7(2)='0' ELSE NOT(OUT_MUX_7);
PP7(12) <= SELECTOR_TABLE_6(2); --PREC
PP7(48) <= '1'; PP7(47) <= NOT (SELECTOR_TABLE_7(2));

PP8(48 DOWNTO 16) <= OUT_MUX_8 WHEN SELECTOR_TABLE_8(2)='0' ELSE NOT(OUT_MUX_8);
PP8(14) <= SELECTOR_TABLE_7(2); --PREC
PP8(50) <= '1'; PP8(49) <= NOT (SELECTOR_TABLE_8(2));

PP9(50 DOWNTO 18) <= OUT_MUX_9 WHEN SELECTOR_TABLE_9(2)='0' ELSE NOT(OUT_MUX_9);
PP9(16) <= SELECTOR_TABLE_8(2); --PREC
PP9(52) <= '1'; PP9(51) <= NOT (SELECTOR_TABLE_9(2));

PP10(52 DOWNTO 20) <= OUT_MUX_10 WHEN SELECTOR_TABLE_10(2)='0' ELSE NOT(OUT_MUX_10);
PP10(18) <= SELECTOR_TABLE_9(2); --PREC
PP10(54) <= '1'; PP10(53) <= NOT (SELECTOR_TABLE_10(2));

PP11(54 DOWNTO 22) <= OUT_MUX_11 WHEN SELECTOR_TABLE_11(2)='0' ELSE NOT(OUT_MUX_11);
PP11(20) <= SELECTOR_TABLE_10(2); --PREC
PP11(56) <= '1'; PP11(55) <= NOT (SELECTOR_TABLE_11(2));

PP12(56 DOWNTO 24) <= OUT_MUX_12 WHEN SELECTOR_TABLE_12(2)='0' ELSE NOT(OUT_MUX_12);
PP12(22) <= SELECTOR_TABLE_11(2); --PREC
PP12(58) <= '1'; PP12(57) <= NOT (SELECTOR_TABLE_12(2));

PP13(58 DOWNTO 26) <= OUT_MUX_13 WHEN SELECTOR_TABLE_13(2)='0' ELSE NOT(OUT_MUX_13);
PP13(24) <= SELECTOR_TABLE_12(2); --PREC
--PARTIAL_PRODUCT_13(25) <= CARRY OUT HALF ADDER;
PP13(60) <= '1'; PP13(59) <= NOT (SELECTOR_TABLE_13(2));

PP14(60 DOWNTO 28) <= OUT_MUX_14 WHEN SELECTOR_TABLE_14(2)='0' ELSE NOT(OUT_MUX_14);
PP14(26) <= SELECTOR_TABLE_13(2); --PREC
--PARTIAL_PRODUCT_14(27) <=  CARRY OUT HALF ADDER;
PP14(62) <= '1'; PP14(61) <= NOT (SELECTOR_TABLE_14(2));

PP15(62 DOWNTO 30) <= OUT_MUX_15 WHEN SELECTOR_TABLE_15(2)='0' ELSE NOT(OUT_MUX_15);
PP15(28) <= SELECTOR_TABLE_14(2); --PREC
--PARTIAL_PRODUCT_15(29,26,27) <= CARRY OUT DI DUE HALF ADDER  
PP15(63) <= NOT (SELECTOR_TABLE_15(2));

PP16(63 DOWNTO 32) <= OUT_MUX_16(31 DOWNTO 0);
PP16(30) <= SELECTOR_TABLE_15(2); --PREC
--PARTIAL_PRODUCT_16(31) <= CARRY OUT  FULL ADDER 
--PARTIAL_PRODUCT_16(29 DOWNTO 28) <= CARRY OUT FULL ADDER

--NEW SCRUCTURE OF PARTIAL PRODUCT (TRIANGLE STRUCTURE)
PARTIAL_PRODUCT_0(63 DOWNTO 0) <= PP16(63 DOWNTO 36) & PP0(35 DOWNTO 0);
PARTIAL_PRODUCT_1(63 DOWNTO 0) <= PP15(63 DOWNTO 37) & PP1(36 DOWNTO 0); 
PARTIAL_PRODUCT_2(62 DOWNTO 2) <= PP14(62 DOWNTO 39) & PP2(38 DOWNTO 2);
PARTIAL_PRODUCT_3(60 DOWNTO 4) <= PP13(60 DOWNTO 41) & PP3(40 DOWNTO 4);
PARTIAL_PRODUCT_4(58 DOWNTO 6) <= PP12(58 DOWNTO 43) & PP4(42 DOWNTO 6);
PARTIAL_PRODUCT_5 (56 DOWNTO 8) <= PP11(56 DOWNTO 45) & PP5(44 DOWNTO 8);
PARTIAL_PRODUCT_6 (54 DOWNTO 10) <= PP10(54 DOWNTO 47) & PP6(46 DOWNTO 10);
PARTIAL_PRODUCT_7 (52 DOWNTO 12) <= PP9(52 DOWNTO 49) & PP7(48 DOWNTO 12);
PARTIAL_PRODUCT_8 (50 DOWNTO 14) <= PP8 (50 DOWNTO 14);
PARTIAL_PRODUCT_9 (48 DOWNTO 16) <= PP9 (48 DOWNTO 16);
PARTIAL_PRODUCT_10 (46 DOWNTO 18) <= PP10 (46 DOWNTO 18);
PARTIAL_PRODUCT_11 (44 DOWNTO 20) <= PP11 (44 DOWNTO 20);
PARTIAL_PRODUCT_12 (42 DOWNTO 22) <= PP12 (42 DOWNTO 22);
PARTIAL_PRODUCT_13 (40 DOWNTO 24) <= PP13 (40 DOWNTO 24);
PARTIAL_PRODUCT_14 (38 DOWNTO 26) <= PP14 (38 DOWNTO 26);
PARTIAL_PRODUCT_15 (36 DOWNTO 28) <= PP15 (36 DOWNTO 28);
PARTIAL_PRODUCT_16 (35 DOWNTO 30) <= PP16 (35 DOWNTO 30);

--LEVEL 6 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--
HA_12_13_24: HA PORT MAP (PARTIAL_PRODUCT_12(24),PARTIAL_PRODUCT_13(24),PARTIAL_PRODUCT_12_1(24),PARTIAL_PRODUCT_11_1(25));
HA_11_12_25: HA PORT MAP (PARTIAL_PRODUCT_11(25),PARTIAL_PRODUCT_12(25),PARTIAL_PRODUCT_12_1(25),PARTIAL_PRODUCT_10_1(26));
HA_13_14_26: HA PORT MAP (PARTIAL_PRODUCT_13(26),PARTIAL_PRODUCT_14(26),PARTIAL_PRODUCT_11_1(26),PARTIAL_PRODUCT_9_1(27));
FA_10_11_12_26: FA PORT MAP (PARTIAL_PRODUCT_10(26),PARTIAL_PRODUCT_11(26),PARTIAL_PRODUCT_12(26),PARTIAL_PRODUCT_12_1(26),PARTIAL_PRODUCT_10_1(27));
HA_12_13_27: HA PORT MAP (PARTIAL_PRODUCT_12(27),PARTIAL_PRODUCT_13(27),PARTIAL_PRODUCT_11_1(27),PARTIAL_PRODUCT_8_1(28));
FA_9_10_11_27: FA PORT MAP (PARTIAL_PRODUCT_9(27),PARTIAL_PRODUCT_10(27),PARTIAL_PRODUCT_11(27),PARTIAL_PRODUCT_12_1(27),PARTIAL_PRODUCT_9_1(28));
HA_14_15_28: HA PORT MAP (PARTIAL_PRODUCT_14(28),PARTIAL_PRODUCT_15(28),PARTIAL_PRODUCT_10_1(28),PARTIAL_PRODUCT_7_1(29));
FA_11_12_13_28: FA PORT MAP (PARTIAL_PRODUCT_11(28),PARTIAL_PRODUCT_12(28),PARTIAL_PRODUCT_13(28),PARTIAL_PRODUCT_11_1(28),PARTIAL_PRODUCT_8_1(29));
FA_8_9_10_28: FA PORT MAP (PARTIAL_PRODUCT_8(28),PARTIAL_PRODUCT_9(28),PARTIAL_PRODUCT_10(28),PARTIAL_PRODUCT_12_1(28),PARTIAL_PRODUCT_9_1(29));
HA_13_14_29: HA PORT MAP (PARTIAL_PRODUCT_13(29),PARTIAL_PRODUCT_14(29),PARTIAL_PRODUCT_10_1(29),PARTIAL_PRODUCT_6_1(30));
FA_10_11_12_29: FA PORT MAP (PARTIAL_PRODUCT_10(29),PARTIAL_PRODUCT_11(29),PARTIAL_PRODUCT_12(29),PARTIAL_PRODUCT_11_1(29),PARTIAL_PRODUCT_7_1(30));
FA_7_8_9_29: FA PORT MAP (PARTIAL_PRODUCT_7(29),PARTIAL_PRODUCT_8(29),PARTIAL_PRODUCT_9(29),PARTIAL_PRODUCT_12_1(29),PARTIAL_PRODUCT_8_1(30));
HA_15_16_30: HA PORT MAP (PARTIAL_PRODUCT_15(30),PARTIAL_PRODUCT_16(30),PARTIAL_PRODUCT_9_1(30),PARTIAL_PRODUCT_5_1(31));
FA_12_13_14_30: FA PORT MAP (PARTIAL_PRODUCT_12(30),PARTIAL_PRODUCT_13(30),PARTIAL_PRODUCT_14(30),PARTIAL_PRODUCT_10_1(30),PARTIAL_PRODUCT_6_1(31));
FA_9_10_11_30: FA PORT MAP (PARTIAL_PRODUCT_9(30),PARTIAL_PRODUCT_10(30),PARTIAL_PRODUCT_11(30),PARTIAL_PRODUCT_11_1(30),PARTIAL_PRODUCT_7_1(31));
FA_6_7_8_30: FA PORT MAP (PARTIAL_PRODUCT_6(30),PARTIAL_PRODUCT_7(30),PARTIAL_PRODUCT_8(30),PARTIAL_PRODUCT_12_1(30),PARTIAL_PRODUCT_8_1(31));
HA_14_15_31: HA PORT MAP (PARTIAL_PRODUCT_14(31),PARTIAL_PRODUCT_15(31),PARTIAL_PRODUCT_9_1(31),PARTIAL_PRODUCT_5_1(32));
FA_11_12_13_31: FA PORT MAP (PARTIAL_PRODUCT_11(31),PARTIAL_PRODUCT_12(31),PARTIAL_PRODUCT_13(31),PARTIAL_PRODUCT_10_1(31),PARTIAL_PRODUCT_6_1(32));
FA_8_9_10_31: FA PORT MAP (PARTIAL_PRODUCT_8(31),PARTIAL_PRODUCT_9(31),PARTIAL_PRODUCT_10(31),PARTIAL_PRODUCT_11_1(31),PARTIAL_PRODUCT_7_1(32));
FA_5_6_7_31: FA PORT MAP (PARTIAL_PRODUCT_5(31),PARTIAL_PRODUCT_6(31),PARTIAL_PRODUCT_7(31),PARTIAL_PRODUCT_12_1(31),PARTIAL_PRODUCT_8_1(32));
FA_14_15_16_32: FA PORT MAP (PARTIAL_PRODUCT_14(32),PARTIAL_PRODUCT_15(32),PARTIAL_PRODUCT_16(32),PARTIAL_PRODUCT_9_1(32),PARTIAL_PRODUCT_5_1(33));
FA_11_12_13_32: FA PORT MAP (PARTIAL_PRODUCT_11(32),PARTIAL_PRODUCT_12(32),PARTIAL_PRODUCT_13(32),PARTIAL_PRODUCT_10_1(32),PARTIAL_PRODUCT_6_1(33));
FA_8_9_10_32: FA PORT MAP (PARTIAL_PRODUCT_8(32),PARTIAL_PRODUCT_9(32),PARTIAL_PRODUCT_10(32),PARTIAL_PRODUCT_11_1(32),PARTIAL_PRODUCT_7_1(33));
FA_5_6_7_32: FA PORT MAP (PARTIAL_PRODUCT_5(32),PARTIAL_PRODUCT_6(32),PARTIAL_PRODUCT_7(32),PARTIAL_PRODUCT_12_1(32),PARTIAL_PRODUCT_8_1(33));
FA_14_15_16_33: FA PORT MAP (PARTIAL_PRODUCT_14(33),PARTIAL_PRODUCT_15(33),PARTIAL_PRODUCT_16(33),PARTIAL_PRODUCT_9_1(33),PARTIAL_PRODUCT_5_1(34));
FA_11_12_13_33: FA PORT MAP (PARTIAL_PRODUCT_11(33),PARTIAL_PRODUCT_12(33),PARTIAL_PRODUCT_13(33),PARTIAL_PRODUCT_10_1(33),PARTIAL_PRODUCT_6_1(34));
FA_8_9_10_33: FA PORT MAP (PARTIAL_PRODUCT_8(33),PARTIAL_PRODUCT_9(33),PARTIAL_PRODUCT_10(33),PARTIAL_PRODUCT_11_1(33),PARTIAL_PRODUCT_7_1(34));
FA_5_6_7_33: FA PORT MAP (PARTIAL_PRODUCT_5(33),PARTIAL_PRODUCT_6(33),PARTIAL_PRODUCT_7(33),PARTIAL_PRODUCT_12_1(33),PARTIAL_PRODUCT_8_1(34));
FA_14_15_16_34: FA PORT MAP (PARTIAL_PRODUCT_14(34),PARTIAL_PRODUCT_15(34),PARTIAL_PRODUCT_16(34),PARTIAL_PRODUCT_9_1(34),PARTIAL_PRODUCT_5_1(35));
FA_11_12_13_34: FA PORT MAP (PARTIAL_PRODUCT_11(34),PARTIAL_PRODUCT_12(34),PARTIAL_PRODUCT_13(34),PARTIAL_PRODUCT_10_1(34),PARTIAL_PRODUCT_6_1(35));
FA_8_9_10_34: FA PORT MAP (PARTIAL_PRODUCT_8(34),PARTIAL_PRODUCT_9(34),PARTIAL_PRODUCT_10(34),PARTIAL_PRODUCT_11_1(34),PARTIAL_PRODUCT_7_1(35));
FA_5_6_7_34: FA PORT MAP (PARTIAL_PRODUCT_5(34),PARTIAL_PRODUCT_6(34),PARTIAL_PRODUCT_7(34),PARTIAL_PRODUCT_12_1(34),PARTIAL_PRODUCT_8_1(35));
FA_14_15_16_35: FA PORT MAP (PARTIAL_PRODUCT_14(35),PARTIAL_PRODUCT_15(35),PARTIAL_PRODUCT_16(35),PARTIAL_PRODUCT_9_1(35),PARTIAL_PRODUCT_5_1(36));
FA_11_12_13_35: FA PORT MAP (PARTIAL_PRODUCT_11(35),PARTIAL_PRODUCT_12(35),PARTIAL_PRODUCT_13(35),PARTIAL_PRODUCT_10_1(35),PARTIAL_PRODUCT_6_1(36));
FA_8_9_10_35: FA PORT MAP (PARTIAL_PRODUCT_8(35),PARTIAL_PRODUCT_9(35),PARTIAL_PRODUCT_10(35),PARTIAL_PRODUCT_11_1(35),PARTIAL_PRODUCT_7_1(36));
FA_5_6_7_35: FA PORT MAP (PARTIAL_PRODUCT_5(35),PARTIAL_PRODUCT_6(35),PARTIAL_PRODUCT_7(35),PARTIAL_PRODUCT_12_1(35),PARTIAL_PRODUCT_8_1(36));
HA_14_15_36: HA PORT MAP (PARTIAL_PRODUCT_14(36),PARTIAL_PRODUCT_15(36),PARTIAL_PRODUCT_9_1(36),PARTIAL_PRODUCT_6_1(37));
FA_11_12_13_36: FA PORT MAP (PARTIAL_PRODUCT_11(36),PARTIAL_PRODUCT_12(36),PARTIAL_PRODUCT_13(36),PARTIAL_PRODUCT_10_1(36),PARTIAL_PRODUCT_7_1(37));
FA_8_9_10_36: FA PORT MAP (PARTIAL_PRODUCT_8(36),PARTIAL_PRODUCT_9(36),PARTIAL_PRODUCT_10(36),PARTIAL_PRODUCT_11_1(36),PARTIAL_PRODUCT_8_1(37));
FA_5_6_7_36: FA PORT MAP (PARTIAL_PRODUCT_5(36),PARTIAL_PRODUCT_6(36),PARTIAL_PRODUCT_7(36),PARTIAL_PRODUCT_12_1(36),PARTIAL_PRODUCT_9_1(37));
FA_12_13_14_37: FA PORT MAP (PARTIAL_PRODUCT_12(37),PARTIAL_PRODUCT_13(37),PARTIAL_PRODUCT_14(37),PARTIAL_PRODUCT_10_1(37),PARTIAL_PRODUCT_7_1(38));
FA_9_10_11_37: FA PORT MAP (PARTIAL_PRODUCT_9(37),PARTIAL_PRODUCT_10(37),PARTIAL_PRODUCT_11(37),PARTIAL_PRODUCT_11_1(37),PARTIAL_PRODUCT_8_1(38));
FA_6_7_8_37: FA PORT MAP (PARTIAL_PRODUCT_6(37),PARTIAL_PRODUCT_7(37),PARTIAL_PRODUCT_8(37),PARTIAL_PRODUCT_12_1(37),PARTIAL_PRODUCT_9_1(38));
HA_13_14_38: HA PORT MAP (PARTIAL_PRODUCT_13(38),PARTIAL_PRODUCT_14(38),PARTIAL_PRODUCT_10_1(38),PARTIAL_PRODUCT_8_1(39));
FA_10_11_12_38: FA PORT MAP (PARTIAL_PRODUCT_10(38),PARTIAL_PRODUCT_11(38),PARTIAL_PRODUCT_12(38),PARTIAL_PRODUCT_11_1(38),PARTIAL_PRODUCT_9_1(39));
FA_7_8_9_38: FA PORT MAP (PARTIAL_PRODUCT_7(38),PARTIAL_PRODUCT_8(38),PARTIAL_PRODUCT_9(38),PARTIAL_PRODUCT_12_1(38),PARTIAL_PRODUCT_10_1(39));
FA_11_12_13_39: FA PORT MAP (PARTIAL_PRODUCT_11(39),PARTIAL_PRODUCT_12(39),PARTIAL_PRODUCT_13(39),PARTIAL_PRODUCT_11_1(39),PARTIAL_PRODUCT_9_1(40));
FA_8_9_10_39: FA PORT MAP (PARTIAL_PRODUCT_8(39),PARTIAL_PRODUCT_9(39),PARTIAL_PRODUCT_10(39),PARTIAL_PRODUCT_12_1(39),PARTIAL_PRODUCT_10_1(40));
HA_12_13_40: HA PORT MAP (PARTIAL_PRODUCT_12(40),PARTIAL_PRODUCT_13(40),PARTIAL_PRODUCT_11_1(40),PARTIAL_PRODUCT_10_1(41));
FA_9_10_11_40: FA PORT MAP (PARTIAL_PRODUCT_9(40),PARTIAL_PRODUCT_10(40),PARTIAL_PRODUCT_11(40),PARTIAL_PRODUCT_12_1(40),PARTIAL_PRODUCT_11_1(41));
FA_10_11_12_41: FA PORT MAP (PARTIAL_PRODUCT_10(41),PARTIAL_PRODUCT_11(41),PARTIAL_PRODUCT_12(41),PARTIAL_PRODUCT_12_1(41),PARTIAL_PRODUCT_11_1(42));
HA_11_12_42: HA PORT MAP (PARTIAL_PRODUCT_11(42),PARTIAL_PRODUCT_12(42),PARTIAL_PRODUCT_12_1(42),PARTIAL_PRODUCT_12_1(43));



PARTIAL_PRODUCT_0_1( 63 downto 0) <= PARTIAL_PRODUCT_0(63 downto 0);
PARTIAL_PRODUCT_1_1( 63 downto 0) <= PARTIAL_PRODUCT_1(63 downto 0); 
PARTIAL_PRODUCT_2_1( 63 downto 0) <= PARTIAL_PRODUCT_2(63 downto 0);
PARTIAL_PRODUCT_3_1( 63 downto 0) <= PARTIAL_PRODUCT_3(63 downto 0);
PARTIAL_PRODUCT_4_1( 63 downto 0) <= PARTIAL_PRODUCT_4(63 downto 0);
PARTIAL_PRODUCT_5_1( 30 downto 0) <= PARTIAL_PRODUCT_5(30 downto 0);
PARTIAL_PRODUCT_6_1( 29 downto 0) <= PARTIAL_PRODUCT_6(29 downto 0); 
PARTIAL_PRODUCT_7_1( 28 downto 0) <= PARTIAL_PRODUCT_7(28 downto 0); 
PARTIAL_PRODUCT_8_1( 27 downto 0) <= PARTIAL_PRODUCT_8(27 downto 0); 
PARTIAL_PRODUCT_9_1( 26 downto 0) <= PARTIAL_PRODUCT_9(26 downto 0); 
PARTIAL_PRODUCT_10_1( 25 downto 0) <= PARTIAL_PRODUCT_10(25 downto 0); 
PARTIAL_PRODUCT_11_1( 24 downto 0) <= PARTIAL_PRODUCT_11(24 downto 0); 
PARTIAL_PRODUCT_12_1( 23 downto 0) <= PARTIAL_PRODUCT_12(23 downto 0); 
PARTIAL_PRODUCT_5_1( 63 downto 37) <= PARTIAL_PRODUCT_5(63 downto 37); 
PARTIAL_PRODUCT_6_1( 63 downto 38) <= PARTIAL_PRODUCT_6(63 downto 38); 
PARTIAL_PRODUCT_7_1( 63 downto 39) <= PARTIAL_PRODUCT_7(63 downto 39); 
PARTIAL_PRODUCT_8_1( 63 downto 40) <= PARTIAL_PRODUCT_8(63 downto 40); 
PARTIAL_PRODUCT_9_1( 63 downto 41) <= PARTIAL_PRODUCT_9(63 downto 41); 
PARTIAL_PRODUCT_10_1( 63 downto 42) <= PARTIAL_PRODUCT_10(63 downto 42); 
PARTIAL_PRODUCT_11_1( 63 downto 43) <= PARTIAL_PRODUCT_11(63 downto 43); 
PARTIAL_PRODUCT_12_1( 63 downto 44) <= PARTIAL_PRODUCT_12(63 downto 44); 

HA_8_9_16_2: HA PORT MAP (PARTIAL_PRODUCT_8_1(16),PARTIAL_PRODUCT_9_1(16),PARTIAL_PRODUCT_8_2(16),PARTIAL_PRODUCT_7_2(17));
HA_7_8_17_2: HA PORT MAP (PARTIAL_PRODUCT_7_1(17),PARTIAL_PRODUCT_8_1(17),PARTIAL_PRODUCT_8_2(17),PARTIAL_PRODUCT_6_2(18));
HA_9_10_18_2: HA PORT MAP (PARTIAL_PRODUCT_9_1(18),PARTIAL_PRODUCT_10_1(18),PARTIAL_PRODUCT_7_2(18),PARTIAL_PRODUCT_5_2(19));
FA_6_7_8_18_2: FA PORT MAP (PARTIAL_PRODUCT_6_1(18),PARTIAL_PRODUCT_7_1(18),PARTIAL_PRODUCT_8_1(18),PARTIAL_PRODUCT_8_2(18),PARTIAL_PRODUCT_6_2(19));
HA_8_9_19_2: HA PORT MAP (PARTIAL_PRODUCT_8_1(19),PARTIAL_PRODUCT_9_1(19),PARTIAL_PRODUCT_7_2(19),PARTIAL_PRODUCT_4_2(20));
FA_5_6_7_19_2: FA PORT MAP (PARTIAL_PRODUCT_5_1(19),PARTIAL_PRODUCT_6_1(19),PARTIAL_PRODUCT_7_1(19),PARTIAL_PRODUCT_8_2(19),PARTIAL_PRODUCT_5_2(20));
HA_10_11_20_2: HA PORT MAP (PARTIAL_PRODUCT_10_1(20),PARTIAL_PRODUCT_11_1(20),PARTIAL_PRODUCT_6_2(20),PARTIAL_PRODUCT_3_2(21));
FA_7_8_9_20_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(20),PARTIAL_PRODUCT_8_1(20),PARTIAL_PRODUCT_9_1(20),PARTIAL_PRODUCT_7_2(20),PARTIAL_PRODUCT_4_2(21));
FA_4_5_6_20_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(20),PARTIAL_PRODUCT_5_1(20),PARTIAL_PRODUCT_6_1(20),PARTIAL_PRODUCT_8_2(20),PARTIAL_PRODUCT_5_2(21));
HA_9_10_21_2: HA PORT MAP (PARTIAL_PRODUCT_9_1(21),PARTIAL_PRODUCT_10_1(21),PARTIAL_PRODUCT_6_2(21),PARTIAL_PRODUCT_2_2(22));
FA_6_7_8_21_2: FA PORT MAP (PARTIAL_PRODUCT_6_1(21),PARTIAL_PRODUCT_7_1(21),PARTIAL_PRODUCT_8_1(21),PARTIAL_PRODUCT_7_2(21),PARTIAL_PRODUCT_3_2(22));
FA_3_4_5_21_2: FA PORT MAP (PARTIAL_PRODUCT_3_1(21),PARTIAL_PRODUCT_4_1(21),PARTIAL_PRODUCT_5_1(21),PARTIAL_PRODUCT_8_2(21),PARTIAL_PRODUCT_4_2(22));
HA_11_12_22_2: HA PORT MAP (PARTIAL_PRODUCT_11_1(22),PARTIAL_PRODUCT_12_1(22),PARTIAL_PRODUCT_5_2(22),PARTIAL_PRODUCT_1_2(23));
FA_8_9_10_22_2: FA PORT MAP (PARTIAL_PRODUCT_8_1(22),PARTIAL_PRODUCT_9_1(22),PARTIAL_PRODUCT_10_1(22),PARTIAL_PRODUCT_6_2(22),PARTIAL_PRODUCT_2_2(23));
FA_5_6_7_22_2: FA PORT MAP (PARTIAL_PRODUCT_5_1(22),PARTIAL_PRODUCT_6_1(22),PARTIAL_PRODUCT_7_1(22),PARTIAL_PRODUCT_7_2(22),PARTIAL_PRODUCT_3_2(23));
FA_2_3_4_22_2: FA PORT MAP (PARTIAL_PRODUCT_2_1(22),PARTIAL_PRODUCT_3_1(22),PARTIAL_PRODUCT_4_1(22),PARTIAL_PRODUCT_8_2(22),PARTIAL_PRODUCT_4_2(23));
HA_10_11_23_2: HA PORT MAP (PARTIAL_PRODUCT_10_1(23),PARTIAL_PRODUCT_11_1(23),PARTIAL_PRODUCT_5_2(23),PARTIAL_PRODUCT_1_2(24));
FA_7_8_9_23_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(23),PARTIAL_PRODUCT_8_1(23),PARTIAL_PRODUCT_9_1(23),PARTIAL_PRODUCT_6_2(23),PARTIAL_PRODUCT_2_2(24));
FA_4_5_6_23_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(23),PARTIAL_PRODUCT_5_1(23),PARTIAL_PRODUCT_6_1(23),PARTIAL_PRODUCT_7_2(23),PARTIAL_PRODUCT_3_2(24));
FA_1_2_3_23_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(23),PARTIAL_PRODUCT_2_1(23),PARTIAL_PRODUCT_3_1(23),PARTIAL_PRODUCT_8_2(23),PARTIAL_PRODUCT_4_2(24));
FA_10_11_12_24_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(24),PARTIAL_PRODUCT_11_1(24),PARTIAL_PRODUCT_12_1(24),PARTIAL_PRODUCT_5_2(24),PARTIAL_PRODUCT_1_2(25));
FA_7_8_9_24_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(24),PARTIAL_PRODUCT_8_1(24),PARTIAL_PRODUCT_9_1(24),PARTIAL_PRODUCT_6_2(24),PARTIAL_PRODUCT_2_2(25));
FA_4_5_6_24_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(24),PARTIAL_PRODUCT_5_1(24),PARTIAL_PRODUCT_6_1(24),PARTIAL_PRODUCT_7_2(24),PARTIAL_PRODUCT_3_2(25));
FA_1_2_3_24_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(24),PARTIAL_PRODUCT_2_1(24),PARTIAL_PRODUCT_3_1(24),PARTIAL_PRODUCT_8_2(24),PARTIAL_PRODUCT_4_2(25));
FA_10_11_12_25_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(25),PARTIAL_PRODUCT_11_1(25),PARTIAL_PRODUCT_12_1(25),PARTIAL_PRODUCT_5_2(25),PARTIAL_PRODUCT_1_2(26));
FA_7_8_9_25_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(25),PARTIAL_PRODUCT_8_1(25),PARTIAL_PRODUCT_9_1(25),PARTIAL_PRODUCT_6_2(25),PARTIAL_PRODUCT_2_2(26));
FA_4_5_6_25_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(25),PARTIAL_PRODUCT_5_1(25),PARTIAL_PRODUCT_6_1(25),PARTIAL_PRODUCT_7_2(25),PARTIAL_PRODUCT_3_2(26));
FA_1_2_3_25_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(25),PARTIAL_PRODUCT_2_1(25),PARTIAL_PRODUCT_3_1(25),PARTIAL_PRODUCT_8_2(25),PARTIAL_PRODUCT_4_2(26));
FA_10_11_12_26_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(26),PARTIAL_PRODUCT_11_1(26),PARTIAL_PRODUCT_12_1(26),PARTIAL_PRODUCT_5_2(26),PARTIAL_PRODUCT_1_2(27));
FA_7_8_9_26_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(26),PARTIAL_PRODUCT_8_1(26),PARTIAL_PRODUCT_9_1(26),PARTIAL_PRODUCT_6_2(26),PARTIAL_PRODUCT_2_2(27));
FA_4_5_6_26_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(26),PARTIAL_PRODUCT_5_1(26),PARTIAL_PRODUCT_6_1(26),PARTIAL_PRODUCT_7_2(26),PARTIAL_PRODUCT_3_2(27));
FA_1_2_3_26_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(26),PARTIAL_PRODUCT_2_1(26),PARTIAL_PRODUCT_3_1(26),PARTIAL_PRODUCT_8_2(26),PARTIAL_PRODUCT_4_2(27));
FA_10_11_12_27_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(27),PARTIAL_PRODUCT_11_1(27),PARTIAL_PRODUCT_12_1(27),PARTIAL_PRODUCT_5_2(27),PARTIAL_PRODUCT_1_2(28));
FA_7_8_9_27_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(27),PARTIAL_PRODUCT_8_1(27),PARTIAL_PRODUCT_9_1(27),PARTIAL_PRODUCT_6_2(27),PARTIAL_PRODUCT_2_2(28));
FA_4_5_6_27_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(27),PARTIAL_PRODUCT_5_1(27),PARTIAL_PRODUCT_6_1(27),PARTIAL_PRODUCT_7_2(27),PARTIAL_PRODUCT_3_2(28));
FA_1_2_3_27_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(27),PARTIAL_PRODUCT_2_1(27),PARTIAL_PRODUCT_3_1(27),PARTIAL_PRODUCT_8_2(27),PARTIAL_PRODUCT_4_2(28));
FA_10_11_12_28_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(28),PARTIAL_PRODUCT_11_1(28),PARTIAL_PRODUCT_12_1(28),PARTIAL_PRODUCT_5_2(28),PARTIAL_PRODUCT_1_2(29));
FA_7_8_9_28_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(28),PARTIAL_PRODUCT_8_1(28),PARTIAL_PRODUCT_9_1(28),PARTIAL_PRODUCT_6_2(28),PARTIAL_PRODUCT_2_2(29));
FA_4_5_6_28_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(28),PARTIAL_PRODUCT_5_1(28),PARTIAL_PRODUCT_6_1(28),PARTIAL_PRODUCT_7_2(28),PARTIAL_PRODUCT_3_2(29));
FA_1_2_3_28_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(28),PARTIAL_PRODUCT_2_1(28),PARTIAL_PRODUCT_3_1(28),PARTIAL_PRODUCT_8_2(28),PARTIAL_PRODUCT_4_2(29));
FA_10_11_12_29_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(29),PARTIAL_PRODUCT_11_1(29),PARTIAL_PRODUCT_12_1(29),PARTIAL_PRODUCT_5_2(29),PARTIAL_PRODUCT_1_2(30));
FA_7_8_9_29_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(29),PARTIAL_PRODUCT_8_1(29),PARTIAL_PRODUCT_9_1(29),PARTIAL_PRODUCT_6_2(29),PARTIAL_PRODUCT_2_2(30));
FA_4_5_6_29_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(29),PARTIAL_PRODUCT_5_1(29),PARTIAL_PRODUCT_6_1(29),PARTIAL_PRODUCT_7_2(29),PARTIAL_PRODUCT_3_2(30));
FA_1_2_3_29_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(29),PARTIAL_PRODUCT_2_1(29),PARTIAL_PRODUCT_3_1(29),PARTIAL_PRODUCT_8_2(29),PARTIAL_PRODUCT_4_2(30));
FA_10_11_12_30_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(30),PARTIAL_PRODUCT_11_1(30),PARTIAL_PRODUCT_12_1(30),PARTIAL_PRODUCT_5_2(30),PARTIAL_PRODUCT_1_2(31));
FA_7_8_9_30_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(30),PARTIAL_PRODUCT_8_1(30),PARTIAL_PRODUCT_9_1(30),PARTIAL_PRODUCT_6_2(30),PARTIAL_PRODUCT_2_2(31));
FA_4_5_6_30_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(30),PARTIAL_PRODUCT_5_1(30),PARTIAL_PRODUCT_6_1(30),PARTIAL_PRODUCT_7_2(30),PARTIAL_PRODUCT_3_2(31));
FA_1_2_3_30_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(30),PARTIAL_PRODUCT_2_1(30),PARTIAL_PRODUCT_3_1(30),PARTIAL_PRODUCT_8_2(30),PARTIAL_PRODUCT_4_2(31));
FA_10_11_12_31_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(31),PARTIAL_PRODUCT_11_1(31),PARTIAL_PRODUCT_12_1(31),PARTIAL_PRODUCT_5_2(31),PARTIAL_PRODUCT_1_2(32));
FA_7_8_9_31_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(31),PARTIAL_PRODUCT_8_1(31),PARTIAL_PRODUCT_9_1(31),PARTIAL_PRODUCT_6_2(31),PARTIAL_PRODUCT_2_2(32));
FA_4_5_6_31_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(31),PARTIAL_PRODUCT_5_1(31),PARTIAL_PRODUCT_6_1(31),PARTIAL_PRODUCT_7_2(31),PARTIAL_PRODUCT_3_2(32));
FA_1_2_3_31_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(31),PARTIAL_PRODUCT_2_1(31),PARTIAL_PRODUCT_3_1(31),PARTIAL_PRODUCT_8_2(31),PARTIAL_PRODUCT_4_2(32));
FA_10_11_12_32_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(32),PARTIAL_PRODUCT_11_1(32),PARTIAL_PRODUCT_12_1(32),PARTIAL_PRODUCT_5_2(32),PARTIAL_PRODUCT_1_2(33));
FA_7_8_9_32_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(32),PARTIAL_PRODUCT_8_1(32),PARTIAL_PRODUCT_9_1(32),PARTIAL_PRODUCT_6_2(32),PARTIAL_PRODUCT_2_2(33));
FA_4_5_6_32_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(32),PARTIAL_PRODUCT_5_1(32),PARTIAL_PRODUCT_6_1(32),PARTIAL_PRODUCT_7_2(32),PARTIAL_PRODUCT_3_2(33));
FA_1_2_3_32_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(32),PARTIAL_PRODUCT_2_1(32),PARTIAL_PRODUCT_3_1(32),PARTIAL_PRODUCT_8_2(32),PARTIAL_PRODUCT_4_2(33));
FA_10_11_12_33_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(33),PARTIAL_PRODUCT_11_1(33),PARTIAL_PRODUCT_12_1(33),PARTIAL_PRODUCT_5_2(33),PARTIAL_PRODUCT_1_2(34));
FA_7_8_9_33_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(33),PARTIAL_PRODUCT_8_1(33),PARTIAL_PRODUCT_9_1(33),PARTIAL_PRODUCT_6_2(33),PARTIAL_PRODUCT_2_2(34));
FA_4_5_6_33_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(33),PARTIAL_PRODUCT_5_1(33),PARTIAL_PRODUCT_6_1(33),PARTIAL_PRODUCT_7_2(33),PARTIAL_PRODUCT_3_2(34));
FA_1_2_3_33_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(33),PARTIAL_PRODUCT_2_1(33),PARTIAL_PRODUCT_3_1(33),PARTIAL_PRODUCT_8_2(33),PARTIAL_PRODUCT_4_2(34));
FA_10_11_12_34_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(34),PARTIAL_PRODUCT_11_1(34),PARTIAL_PRODUCT_12_1(34),PARTIAL_PRODUCT_5_2(34),PARTIAL_PRODUCT_1_2(35));
FA_7_8_9_34_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(34),PARTIAL_PRODUCT_8_1(34),PARTIAL_PRODUCT_9_1(34),PARTIAL_PRODUCT_6_2(34),PARTIAL_PRODUCT_2_2(35));
FA_4_5_6_34_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(34),PARTIAL_PRODUCT_5_1(34),PARTIAL_PRODUCT_6_1(34),PARTIAL_PRODUCT_7_2(34),PARTIAL_PRODUCT_3_2(35));
FA_1_2_3_34_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(34),PARTIAL_PRODUCT_2_1(34),PARTIAL_PRODUCT_3_1(34),PARTIAL_PRODUCT_8_2(34),PARTIAL_PRODUCT_4_2(35));
FA_10_11_12_35_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(35),PARTIAL_PRODUCT_11_1(35),PARTIAL_PRODUCT_12_1(35),PARTIAL_PRODUCT_5_2(35),PARTIAL_PRODUCT_1_2(36));
FA_7_8_9_35_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(35),PARTIAL_PRODUCT_8_1(35),PARTIAL_PRODUCT_9_1(35),PARTIAL_PRODUCT_6_2(35),PARTIAL_PRODUCT_2_2(36));
FA_4_5_6_35_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(35),PARTIAL_PRODUCT_5_1(35),PARTIAL_PRODUCT_6_1(35),PARTIAL_PRODUCT_7_2(35),PARTIAL_PRODUCT_3_2(36));
FA_1_2_3_35_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(35),PARTIAL_PRODUCT_2_1(35),PARTIAL_PRODUCT_3_1(35),PARTIAL_PRODUCT_8_2(35),PARTIAL_PRODUCT_4_2(36));
FA_10_11_12_36_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(36),PARTIAL_PRODUCT_11_1(36),PARTIAL_PRODUCT_12_1(36),PARTIAL_PRODUCT_5_2(36),PARTIAL_PRODUCT_1_2(37));
FA_7_8_9_36_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(36),PARTIAL_PRODUCT_8_1(36),PARTIAL_PRODUCT_9_1(36),PARTIAL_PRODUCT_6_2(36),PARTIAL_PRODUCT_2_2(37));
FA_4_5_6_36_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(36),PARTIAL_PRODUCT_5_1(36),PARTIAL_PRODUCT_6_1(36),PARTIAL_PRODUCT_7_2(36),PARTIAL_PRODUCT_3_2(37));
FA_1_2_3_36_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(36),PARTIAL_PRODUCT_2_1(36),PARTIAL_PRODUCT_3_1(36),PARTIAL_PRODUCT_8_2(36),PARTIAL_PRODUCT_4_2(37));
FA_10_11_12_37_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(37),PARTIAL_PRODUCT_11_1(37),PARTIAL_PRODUCT_12_1(37),PARTIAL_PRODUCT_5_2(37),PARTIAL_PRODUCT_1_2(38));
FA_7_8_9_37_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(37),PARTIAL_PRODUCT_8_1(37),PARTIAL_PRODUCT_9_1(37),PARTIAL_PRODUCT_6_2(37),PARTIAL_PRODUCT_2_2(38));
FA_4_5_6_37_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(37),PARTIAL_PRODUCT_5_1(37),PARTIAL_PRODUCT_6_1(37),PARTIAL_PRODUCT_7_2(37),PARTIAL_PRODUCT_3_2(38));
FA_1_2_3_37_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(37),PARTIAL_PRODUCT_2_1(37),PARTIAL_PRODUCT_3_1(37),PARTIAL_PRODUCT_8_2(37),PARTIAL_PRODUCT_4_2(38));
FA_10_11_12_38_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(38),PARTIAL_PRODUCT_11_1(38),PARTIAL_PRODUCT_12_1(38),PARTIAL_PRODUCT_5_2(38),PARTIAL_PRODUCT_1_2(39));
FA_7_8_9_38_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(38),PARTIAL_PRODUCT_8_1(38),PARTIAL_PRODUCT_9_1(38),PARTIAL_PRODUCT_6_2(38),PARTIAL_PRODUCT_2_2(39));
FA_4_5_6_38_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(38),PARTIAL_PRODUCT_5_1(38),PARTIAL_PRODUCT_6_1(38),PARTIAL_PRODUCT_7_2(38),PARTIAL_PRODUCT_3_2(39));
FA_1_2_3_38_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(38),PARTIAL_PRODUCT_2_1(38),PARTIAL_PRODUCT_3_1(38),PARTIAL_PRODUCT_8_2(38),PARTIAL_PRODUCT_4_2(39));
FA_10_11_12_39_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(39),PARTIAL_PRODUCT_11_1(39),PARTIAL_PRODUCT_12_1(39),PARTIAL_PRODUCT_5_2(39),PARTIAL_PRODUCT_1_2(40));
FA_7_8_9_39_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(39),PARTIAL_PRODUCT_8_1(39),PARTIAL_PRODUCT_9_1(39),PARTIAL_PRODUCT_6_2(39),PARTIAL_PRODUCT_2_2(40));
FA_4_5_6_39_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(39),PARTIAL_PRODUCT_5_1(39),PARTIAL_PRODUCT_6_1(39),PARTIAL_PRODUCT_7_2(39),PARTIAL_PRODUCT_3_2(40));
FA_1_2_3_39_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(39),PARTIAL_PRODUCT_2_1(39),PARTIAL_PRODUCT_3_1(39),PARTIAL_PRODUCT_8_2(39),PARTIAL_PRODUCT_4_2(40));
FA_10_11_12_40_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(40),PARTIAL_PRODUCT_11_1(40),PARTIAL_PRODUCT_12_1(40),PARTIAL_PRODUCT_5_2(40),PARTIAL_PRODUCT_1_2(41));
FA_7_8_9_40_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(40),PARTIAL_PRODUCT_8_1(40),PARTIAL_PRODUCT_9_1(40),PARTIAL_PRODUCT_6_2(40),PARTIAL_PRODUCT_2_2(41));
FA_4_5_6_40_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(40),PARTIAL_PRODUCT_5_1(40),PARTIAL_PRODUCT_6_1(40),PARTIAL_PRODUCT_7_2(40),PARTIAL_PRODUCT_3_2(41));
FA_1_2_3_40_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(40),PARTIAL_PRODUCT_2_1(40),PARTIAL_PRODUCT_3_1(40),PARTIAL_PRODUCT_8_2(40),PARTIAL_PRODUCT_4_2(41));
FA_10_11_12_41_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(41),PARTIAL_PRODUCT_11_1(41),PARTIAL_PRODUCT_12_1(41),PARTIAL_PRODUCT_5_2(41),PARTIAL_PRODUCT_1_2(42));
FA_7_8_9_41_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(41),PARTIAL_PRODUCT_8_1(41),PARTIAL_PRODUCT_9_1(41),PARTIAL_PRODUCT_6_2(41),PARTIAL_PRODUCT_2_2(42));
FA_4_5_6_41_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(41),PARTIAL_PRODUCT_5_1(41),PARTIAL_PRODUCT_6_1(41),PARTIAL_PRODUCT_7_2(41),PARTIAL_PRODUCT_3_2(42));
FA_1_2_3_41_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(41),PARTIAL_PRODUCT_2_1(41),PARTIAL_PRODUCT_3_1(41),PARTIAL_PRODUCT_8_2(41),PARTIAL_PRODUCT_4_2(42));
FA_10_11_12_42_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(42),PARTIAL_PRODUCT_11_1(42),PARTIAL_PRODUCT_12_1(42),PARTIAL_PRODUCT_5_2(42),PARTIAL_PRODUCT_1_2(43));
FA_7_8_9_42_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(42),PARTIAL_PRODUCT_8_1(42),PARTIAL_PRODUCT_9_1(42),PARTIAL_PRODUCT_6_2(42),PARTIAL_PRODUCT_2_2(43));
FA_4_5_6_42_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(42),PARTIAL_PRODUCT_5_1(42),PARTIAL_PRODUCT_6_1(42),PARTIAL_PRODUCT_7_2(42),PARTIAL_PRODUCT_3_2(43));
FA_1_2_3_42_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(42),PARTIAL_PRODUCT_2_1(42),PARTIAL_PRODUCT_3_1(42),PARTIAL_PRODUCT_8_2(42),PARTIAL_PRODUCT_4_2(43));
FA_10_11_12_43_2: FA PORT MAP (PARTIAL_PRODUCT_10_1(43),PARTIAL_PRODUCT_11_1(43),PARTIAL_PRODUCT_12_1(43),PARTIAL_PRODUCT_5_2(43),PARTIAL_PRODUCT_1_2(44));
FA_7_8_9_43_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(43),PARTIAL_PRODUCT_8_1(43),PARTIAL_PRODUCT_9_1(43),PARTIAL_PRODUCT_6_2(43),PARTIAL_PRODUCT_2_2(44));
FA_4_5_6_43_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(43),PARTIAL_PRODUCT_5_1(43),PARTIAL_PRODUCT_6_1(43),PARTIAL_PRODUCT_7_2(43),PARTIAL_PRODUCT_3_2(44));
FA_1_2_3_43_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(43),PARTIAL_PRODUCT_2_1(43),PARTIAL_PRODUCT_3_1(43),PARTIAL_PRODUCT_8_2(43),PARTIAL_PRODUCT_4_2(44));
HA_10_11_44_2: HA PORT MAP (PARTIAL_PRODUCT_10_1(44),PARTIAL_PRODUCT_11_1(44),PARTIAL_PRODUCT_5_2(44),PARTIAL_PRODUCT_2_2(45));
FA_7_8_9_44_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(44),PARTIAL_PRODUCT_8_1(44),PARTIAL_PRODUCT_9_1(44),PARTIAL_PRODUCT_6_2(44),PARTIAL_PRODUCT_3_2(45));
FA_4_5_6_44_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(44),PARTIAL_PRODUCT_5_1(44),PARTIAL_PRODUCT_6_1(44),PARTIAL_PRODUCT_7_2(44),PARTIAL_PRODUCT_4_2(45));
FA_1_2_3_44_2: FA PORT MAP (PARTIAL_PRODUCT_1_1(44),PARTIAL_PRODUCT_2_1(44),PARTIAL_PRODUCT_3_1(44),PARTIAL_PRODUCT_8_2(44),PARTIAL_PRODUCT_5_2(45));
FA_8_9_10_45_2: FA PORT MAP (PARTIAL_PRODUCT_8_1(45),PARTIAL_PRODUCT_9_1(45),PARTIAL_PRODUCT_10_1(45),PARTIAL_PRODUCT_6_2(45),PARTIAL_PRODUCT_3_2(46));
FA_5_6_7_45_2: FA PORT MAP (PARTIAL_PRODUCT_5_1(45),PARTIAL_PRODUCT_6_1(45),PARTIAL_PRODUCT_7_1(45),PARTIAL_PRODUCT_7_2(45),PARTIAL_PRODUCT_4_2(46));
FA_2_3_4_45_2: FA PORT MAP (PARTIAL_PRODUCT_2_1(45),PARTIAL_PRODUCT_3_1(45),PARTIAL_PRODUCT_4_1(45),PARTIAL_PRODUCT_8_2(45),PARTIAL_PRODUCT_5_2(46));
HA_9_10_46_2: HA PORT MAP (PARTIAL_PRODUCT_9_1(46),PARTIAL_PRODUCT_10_1(46),PARTIAL_PRODUCT_6_2(46),PARTIAL_PRODUCT_4_2(47));
FA_6_7_8_46_2: FA PORT MAP (PARTIAL_PRODUCT_6_1(46),PARTIAL_PRODUCT_7_1(46),PARTIAL_PRODUCT_8_1(46),PARTIAL_PRODUCT_7_2(46),PARTIAL_PRODUCT_5_2(47));
FA_3_4_5_46_2: FA PORT MAP (PARTIAL_PRODUCT_3_1(46),PARTIAL_PRODUCT_4_1(46),PARTIAL_PRODUCT_5_1(46),PARTIAL_PRODUCT_8_2(46),PARTIAL_PRODUCT_6_2(47));
FA_7_8_9_47_2: FA PORT MAP (PARTIAL_PRODUCT_7_1(47),PARTIAL_PRODUCT_8_1(47),PARTIAL_PRODUCT_9_1(47),PARTIAL_PRODUCT_7_2(47),PARTIAL_PRODUCT_5_2(48));
FA_4_5_6_47_2: FA PORT MAP (PARTIAL_PRODUCT_4_1(47),PARTIAL_PRODUCT_5_1(47),PARTIAL_PRODUCT_6_1(47),PARTIAL_PRODUCT_8_2(47),PARTIAL_PRODUCT_6_2(48));
HA_8_9_48_2: HA PORT MAP (PARTIAL_PRODUCT_8_1(48),PARTIAL_PRODUCT_9_1(48),PARTIAL_PRODUCT_7_2(48),PARTIAL_PRODUCT_6_2(49));
FA_5_6_7_48_2: FA PORT MAP (PARTIAL_PRODUCT_5_1(48),PARTIAL_PRODUCT_6_1(48),PARTIAL_PRODUCT_7_1(48),PARTIAL_PRODUCT_8_2(48),PARTIAL_PRODUCT_7_2(49));
FA_6_7_8_49_2: FA PORT MAP (PARTIAL_PRODUCT_6_1(49),PARTIAL_PRODUCT_7_1(49),PARTIAL_PRODUCT_8_1(49),PARTIAL_PRODUCT_8_2(49),PARTIAL_PRODUCT_7_2(50));
HA_7_8_50_2: HA PORT MAP (PARTIAL_PRODUCT_7_1(50),PARTIAL_PRODUCT_8_1(50),PARTIAL_PRODUCT_8_2(50),PARTIAL_PRODUCT_8_2(51));

PARTIAL_PRODUCT_0_2( 63 downto 0) <= PARTIAL_PRODUCT_0_1(63 downto 0); 
PARTIAL_PRODUCT_1_2( 22 downto 0) <= PARTIAL_PRODUCT_1_1(22 downto 0); 
PARTIAL_PRODUCT_2_2( 21 downto 0) <= PARTIAL_PRODUCT_2_1(21 downto 0); 
PARTIAL_PRODUCT_3_2( 20 downto 0) <= PARTIAL_PRODUCT_3_1(20 downto 0); 
PARTIAL_PRODUCT_4_2( 19 downto 0) <= PARTIAL_PRODUCT_4_1(19 downto 0); 
PARTIAL_PRODUCT_5_2( 18 downto 0) <= PARTIAL_PRODUCT_5_1(18 downto 0); 
PARTIAL_PRODUCT_6_2( 17 downto 0) <= PARTIAL_PRODUCT_6_1(17 downto 0); 
PARTIAL_PRODUCT_7_2( 16 downto 0) <= PARTIAL_PRODUCT_7_1(16 downto 0); 
PARTIAL_PRODUCT_8_2( 15 downto 0) <= PARTIAL_PRODUCT_8_1(15 downto 0); 
PARTIAL_PRODUCT_1_2( 63 downto 45) <= PARTIAL_PRODUCT_1_1(63 downto 45); 
PARTIAL_PRODUCT_2_2( 63 downto 46) <= PARTIAL_PRODUCT_2_1(63 downto 46); 
PARTIAL_PRODUCT_3_2( 63 downto 47) <= PARTIAL_PRODUCT_3_1(63 downto 47); 
PARTIAL_PRODUCT_4_2( 63 downto 48) <= PARTIAL_PRODUCT_4_1(63 downto 48); 
PARTIAL_PRODUCT_5_2( 63 downto 49) <= PARTIAL_PRODUCT_5_1(63 downto 49); 
PARTIAL_PRODUCT_6_2( 63 downto 50) <= PARTIAL_PRODUCT_6_1(63 downto 50); 
PARTIAL_PRODUCT_7_2( 63 downto 51) <= PARTIAL_PRODUCT_7_1(63 downto 51); 
PARTIAL_PRODUCT_8_2( 63 downto 52) <= PARTIAL_PRODUCT_8_1(63 downto 52); 

HA_5_6_10_3: HA PORT MAP (PARTIAL_PRODUCT_5_2(10),PARTIAL_PRODUCT_6_2(10),PARTIAL_PRODUCT_5_3(10),PARTIAL_PRODUCT_4_3(11));
HA_4_5_11_3: HA PORT MAP (PARTIAL_PRODUCT_4_2(11),PARTIAL_PRODUCT_5_2(11),PARTIAL_PRODUCT_5_3(11),PARTIAL_PRODUCT_3_3(12));
HA_6_7_12_3: HA PORT MAP (PARTIAL_PRODUCT_6_2(12),PARTIAL_PRODUCT_7_2(12),PARTIAL_PRODUCT_4_3(12),PARTIAL_PRODUCT_2_3(13));
FA_3_4_5_12_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(12),PARTIAL_PRODUCT_4_2(12),PARTIAL_PRODUCT_5_2(12),PARTIAL_PRODUCT_5_3(12),PARTIAL_PRODUCT_3_3(13));
HA_5_6_13_3: HA PORT MAP (PARTIAL_PRODUCT_5_2(13),PARTIAL_PRODUCT_6_2(13),PARTIAL_PRODUCT_4_3(13),PARTIAL_PRODUCT_1_3(14));
FA_2_3_4_13_3: FA PORT MAP (PARTIAL_PRODUCT_2_2(13),PARTIAL_PRODUCT_3_2(13),PARTIAL_PRODUCT_4_2(13),PARTIAL_PRODUCT_5_3(13),PARTIAL_PRODUCT_2_3(14));
HA_7_8_14_3: HA PORT MAP (PARTIAL_PRODUCT_7_2(14),PARTIAL_PRODUCT_8_2(14),PARTIAL_PRODUCT_3_3(14),PARTIAL_PRODUCT_0_3(15));
FA_4_5_6_14_3: FA PORT MAP (PARTIAL_PRODUCT_4_2(14),PARTIAL_PRODUCT_5_2(14),PARTIAL_PRODUCT_6_2(14),PARTIAL_PRODUCT_4_3(14),PARTIAL_PRODUCT_1_3(15));
FA_1_2_3_14_3: FA PORT MAP (PARTIAL_PRODUCT_1_2(14),PARTIAL_PRODUCT_2_2(14),PARTIAL_PRODUCT_3_2(14),PARTIAL_PRODUCT_5_3(14),PARTIAL_PRODUCT_2_3(15));
HA_6_7_15_3: HA PORT MAP (PARTIAL_PRODUCT_6_2(15),PARTIAL_PRODUCT_7_2(15),PARTIAL_PRODUCT_3_3(15),PARTIAL_PRODUCT_0_3(16));
FA_3_4_5_15_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(15),PARTIAL_PRODUCT_4_2(15),PARTIAL_PRODUCT_5_2(15),PARTIAL_PRODUCT_4_3(15),PARTIAL_PRODUCT_1_3(16));
FA_0_1_2_15_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(15),PARTIAL_PRODUCT_1_2(15),PARTIAL_PRODUCT_2_2(15),PARTIAL_PRODUCT_5_3(15),PARTIAL_PRODUCT_2_3(16));
FA_6_7_8_16_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(16),PARTIAL_PRODUCT_7_2(16),PARTIAL_PRODUCT_8_2(16),PARTIAL_PRODUCT_3_3(16),PARTIAL_PRODUCT_0_3(17));
FA_3_4_5_16_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(16),PARTIAL_PRODUCT_4_2(16),PARTIAL_PRODUCT_5_2(16),PARTIAL_PRODUCT_4_3(16),PARTIAL_PRODUCT_1_3(17));
FA_0_1_2_16_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(16),PARTIAL_PRODUCT_1_2(16),PARTIAL_PRODUCT_2_2(16),PARTIAL_PRODUCT_5_3(16),PARTIAL_PRODUCT_2_3(17));
FA_6_7_8_17_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(17),PARTIAL_PRODUCT_7_2(17),PARTIAL_PRODUCT_8_2(17),PARTIAL_PRODUCT_3_3(17),PARTIAL_PRODUCT_0_3(18));
FA_3_4_5_17_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(17),PARTIAL_PRODUCT_4_2(17),PARTIAL_PRODUCT_5_2(17),PARTIAL_PRODUCT_4_3(17),PARTIAL_PRODUCT_1_3(18));
FA_0_1_2_17_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(17),PARTIAL_PRODUCT_1_2(17),PARTIAL_PRODUCT_2_2(17),PARTIAL_PRODUCT_5_3(17),PARTIAL_PRODUCT_2_3(18));
FA_6_7_8_18_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(18),PARTIAL_PRODUCT_7_2(18),PARTIAL_PRODUCT_8_2(18),PARTIAL_PRODUCT_3_3(18),PARTIAL_PRODUCT_0_3(19));
FA_3_4_5_18_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(18),PARTIAL_PRODUCT_4_2(18),PARTIAL_PRODUCT_5_2(18),PARTIAL_PRODUCT_4_3(18),PARTIAL_PRODUCT_1_3(19));
FA_0_1_2_18_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(18),PARTIAL_PRODUCT_1_2(18),PARTIAL_PRODUCT_2_2(18),PARTIAL_PRODUCT_5_3(18),PARTIAL_PRODUCT_2_3(19));
FA_6_7_8_19_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(19),PARTIAL_PRODUCT_7_2(19),PARTIAL_PRODUCT_8_2(19),PARTIAL_PRODUCT_3_3(19),PARTIAL_PRODUCT_0_3(20));
FA_3_4_5_19_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(19),PARTIAL_PRODUCT_4_2(19),PARTIAL_PRODUCT_5_2(19),PARTIAL_PRODUCT_4_3(19),PARTIAL_PRODUCT_1_3(20));
FA_0_1_2_19_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(19),PARTIAL_PRODUCT_1_2(19),PARTIAL_PRODUCT_2_2(19),PARTIAL_PRODUCT_5_3(19),PARTIAL_PRODUCT_2_3(20));
FA_6_7_8_20_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(20),PARTIAL_PRODUCT_7_2(20),PARTIAL_PRODUCT_8_2(20),PARTIAL_PRODUCT_3_3(20),PARTIAL_PRODUCT_0_3(21));
FA_3_4_5_20_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(20),PARTIAL_PRODUCT_4_2(20),PARTIAL_PRODUCT_5_2(20),PARTIAL_PRODUCT_4_3(20),PARTIAL_PRODUCT_1_3(21));
FA_0_1_2_20_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(20),PARTIAL_PRODUCT_1_2(20),PARTIAL_PRODUCT_2_2(20),PARTIAL_PRODUCT_5_3(20),PARTIAL_PRODUCT_2_3(21));
FA_6_7_8_21_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(21),PARTIAL_PRODUCT_7_2(21),PARTIAL_PRODUCT_8_2(21),PARTIAL_PRODUCT_3_3(21),PARTIAL_PRODUCT_0_3(22));
FA_3_4_5_21_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(21),PARTIAL_PRODUCT_4_2(21),PARTIAL_PRODUCT_5_2(21),PARTIAL_PRODUCT_4_3(21),PARTIAL_PRODUCT_1_3(22));
FA_0_1_2_21_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(21),PARTIAL_PRODUCT_1_2(21),PARTIAL_PRODUCT_2_2(21),PARTIAL_PRODUCT_5_3(21),PARTIAL_PRODUCT_2_3(22));
FA_6_7_8_22_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(22),PARTIAL_PRODUCT_7_2(22),PARTIAL_PRODUCT_8_2(22),PARTIAL_PRODUCT_3_3(22),PARTIAL_PRODUCT_0_3(23));
FA_3_4_5_22_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(22),PARTIAL_PRODUCT_4_2(22),PARTIAL_PRODUCT_5_2(22),PARTIAL_PRODUCT_4_3(22),PARTIAL_PRODUCT_1_3(23));
FA_0_1_2_22_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(22),PARTIAL_PRODUCT_1_2(22),PARTIAL_PRODUCT_2_2(22),PARTIAL_PRODUCT_5_3(22),PARTIAL_PRODUCT_2_3(23));
FA_6_7_8_23_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(23),PARTIAL_PRODUCT_7_2(23),PARTIAL_PRODUCT_8_2(23),PARTIAL_PRODUCT_3_3(23),PARTIAL_PRODUCT_0_3(24));
FA_3_4_5_23_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(23),PARTIAL_PRODUCT_4_2(23),PARTIAL_PRODUCT_5_2(23),PARTIAL_PRODUCT_4_3(23),PARTIAL_PRODUCT_1_3(24));
FA_0_1_2_23_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(23),PARTIAL_PRODUCT_1_2(23),PARTIAL_PRODUCT_2_2(23),PARTIAL_PRODUCT_5_3(23),PARTIAL_PRODUCT_2_3(24));
FA_6_7_8_24_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(24),PARTIAL_PRODUCT_7_2(24),PARTIAL_PRODUCT_8_2(24),PARTIAL_PRODUCT_3_3(24),PARTIAL_PRODUCT_0_3(25));
FA_3_4_5_24_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(24),PARTIAL_PRODUCT_4_2(24),PARTIAL_PRODUCT_5_2(24),PARTIAL_PRODUCT_4_3(24),PARTIAL_PRODUCT_1_3(25));
FA_0_1_2_24_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(24),PARTIAL_PRODUCT_1_2(24),PARTIAL_PRODUCT_2_2(24),PARTIAL_PRODUCT_5_3(24),PARTIAL_PRODUCT_2_3(25));
FA_6_7_8_25_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(25),PARTIAL_PRODUCT_7_2(25),PARTIAL_PRODUCT_8_2(25),PARTIAL_PRODUCT_3_3(25),PARTIAL_PRODUCT_0_3(26));
FA_3_4_5_25_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(25),PARTIAL_PRODUCT_4_2(25),PARTIAL_PRODUCT_5_2(25),PARTIAL_PRODUCT_4_3(25),PARTIAL_PRODUCT_1_3(26));
FA_0_1_2_25_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(25),PARTIAL_PRODUCT_1_2(25),PARTIAL_PRODUCT_2_2(25),PARTIAL_PRODUCT_5_3(25),PARTIAL_PRODUCT_2_3(26));
FA_6_7_8_26_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(26),PARTIAL_PRODUCT_7_2(26),PARTIAL_PRODUCT_8_2(26),PARTIAL_PRODUCT_3_3(26),PARTIAL_PRODUCT_0_3(27));
FA_3_4_5_26_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(26),PARTIAL_PRODUCT_4_2(26),PARTIAL_PRODUCT_5_2(26),PARTIAL_PRODUCT_4_3(26),PARTIAL_PRODUCT_1_3(27));
FA_0_1_2_26_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(26),PARTIAL_PRODUCT_1_2(26),PARTIAL_PRODUCT_2_2(26),PARTIAL_PRODUCT_5_3(26),PARTIAL_PRODUCT_2_3(27));
FA_6_7_8_27_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(27),PARTIAL_PRODUCT_7_2(27),PARTIAL_PRODUCT_8_2(27),PARTIAL_PRODUCT_3_3(27),PARTIAL_PRODUCT_0_3(28));
FA_3_4_5_27_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(27),PARTIAL_PRODUCT_4_2(27),PARTIAL_PRODUCT_5_2(27),PARTIAL_PRODUCT_4_3(27),PARTIAL_PRODUCT_1_3(28));
FA_0_1_2_27_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(27),PARTIAL_PRODUCT_1_2(27),PARTIAL_PRODUCT_2_2(27),PARTIAL_PRODUCT_5_3(27),PARTIAL_PRODUCT_2_3(28));
FA_6_7_8_28_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(28),PARTIAL_PRODUCT_7_2(28),PARTIAL_PRODUCT_8_2(28),PARTIAL_PRODUCT_3_3(28),PARTIAL_PRODUCT_0_3(29));
FA_3_4_5_28_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(28),PARTIAL_PRODUCT_4_2(28),PARTIAL_PRODUCT_5_2(28),PARTIAL_PRODUCT_4_3(28),PARTIAL_PRODUCT_1_3(29));
FA_0_1_2_28_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(28),PARTIAL_PRODUCT_1_2(28),PARTIAL_PRODUCT_2_2(28),PARTIAL_PRODUCT_5_3(28),PARTIAL_PRODUCT_2_3(29));
FA_6_7_8_29_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(29),PARTIAL_PRODUCT_7_2(29),PARTIAL_PRODUCT_8_2(29),PARTIAL_PRODUCT_3_3(29),PARTIAL_PRODUCT_0_3(30));
FA_3_4_5_29_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(29),PARTIAL_PRODUCT_4_2(29),PARTIAL_PRODUCT_5_2(29),PARTIAL_PRODUCT_4_3(29),PARTIAL_PRODUCT_1_3(30));
FA_0_1_2_29_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(29),PARTIAL_PRODUCT_1_2(29),PARTIAL_PRODUCT_2_2(29),PARTIAL_PRODUCT_5_3(29),PARTIAL_PRODUCT_2_3(30));
FA_6_7_8_30_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(30),PARTIAL_PRODUCT_7_2(30),PARTIAL_PRODUCT_8_2(30),PARTIAL_PRODUCT_3_3(30),PARTIAL_PRODUCT_0_3(31));
FA_3_4_5_30_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(30),PARTIAL_PRODUCT_4_2(30),PARTIAL_PRODUCT_5_2(30),PARTIAL_PRODUCT_4_3(30),PARTIAL_PRODUCT_1_3(31));
FA_0_1_2_30_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(30),PARTIAL_PRODUCT_1_2(30),PARTIAL_PRODUCT_2_2(30),PARTIAL_PRODUCT_5_3(30),PARTIAL_PRODUCT_2_3(31));
FA_6_7_8_31_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(31),PARTIAL_PRODUCT_7_2(31),PARTIAL_PRODUCT_8_2(31),PARTIAL_PRODUCT_3_3(31),PARTIAL_PRODUCT_0_3(32));
FA_3_4_5_31_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(31),PARTIAL_PRODUCT_4_2(31),PARTIAL_PRODUCT_5_2(31),PARTIAL_PRODUCT_4_3(31),PARTIAL_PRODUCT_1_3(32));
FA_0_1_2_31_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(31),PARTIAL_PRODUCT_1_2(31),PARTIAL_PRODUCT_2_2(31),PARTIAL_PRODUCT_5_3(31),PARTIAL_PRODUCT_2_3(32));
FA_6_7_8_32_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(32),PARTIAL_PRODUCT_7_2(32),PARTIAL_PRODUCT_8_2(32),PARTIAL_PRODUCT_3_3(32),PARTIAL_PRODUCT_0_3(33));
FA_3_4_5_32_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(32),PARTIAL_PRODUCT_4_2(32),PARTIAL_PRODUCT_5_2(32),PARTIAL_PRODUCT_4_3(32),PARTIAL_PRODUCT_1_3(33));
FA_0_1_2_32_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(32),PARTIAL_PRODUCT_1_2(32),PARTIAL_PRODUCT_2_2(32),PARTIAL_PRODUCT_5_3(32),PARTIAL_PRODUCT_2_3(33));
FA_6_7_8_33_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(33),PARTIAL_PRODUCT_7_2(33),PARTIAL_PRODUCT_8_2(33),PARTIAL_PRODUCT_3_3(33),PARTIAL_PRODUCT_0_3(34));
FA_3_4_5_33_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(33),PARTIAL_PRODUCT_4_2(33),PARTIAL_PRODUCT_5_2(33),PARTIAL_PRODUCT_4_3(33),PARTIAL_PRODUCT_1_3(34));
FA_0_1_2_33_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(33),PARTIAL_PRODUCT_1_2(33),PARTIAL_PRODUCT_2_2(33),PARTIAL_PRODUCT_5_3(33),PARTIAL_PRODUCT_2_3(34));
FA_6_7_8_34_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(34),PARTIAL_PRODUCT_7_2(34),PARTIAL_PRODUCT_8_2(34),PARTIAL_PRODUCT_3_3(34),PARTIAL_PRODUCT_0_3(35));
FA_3_4_5_34_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(34),PARTIAL_PRODUCT_4_2(34),PARTIAL_PRODUCT_5_2(34),PARTIAL_PRODUCT_4_3(34),PARTIAL_PRODUCT_1_3(35));
FA_0_1_2_34_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(34),PARTIAL_PRODUCT_1_2(34),PARTIAL_PRODUCT_2_2(34),PARTIAL_PRODUCT_5_3(34),PARTIAL_PRODUCT_2_3(35));
FA_6_7_8_35_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(35),PARTIAL_PRODUCT_7_2(35),PARTIAL_PRODUCT_8_2(35),PARTIAL_PRODUCT_3_3(35),PARTIAL_PRODUCT_0_3(36));
FA_3_4_5_35_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(35),PARTIAL_PRODUCT_4_2(35),PARTIAL_PRODUCT_5_2(35),PARTIAL_PRODUCT_4_3(35),PARTIAL_PRODUCT_1_3(36));
FA_0_1_2_35_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(35),PARTIAL_PRODUCT_1_2(35),PARTIAL_PRODUCT_2_2(35),PARTIAL_PRODUCT_5_3(35),PARTIAL_PRODUCT_2_3(36));
FA_6_7_8_36_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(36),PARTIAL_PRODUCT_7_2(36),PARTIAL_PRODUCT_8_2(36),PARTIAL_PRODUCT_3_3(36),PARTIAL_PRODUCT_0_3(37));
FA_3_4_5_36_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(36),PARTIAL_PRODUCT_4_2(36),PARTIAL_PRODUCT_5_2(36),PARTIAL_PRODUCT_4_3(36),PARTIAL_PRODUCT_1_3(37));
FA_0_1_2_36_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(36),PARTIAL_PRODUCT_1_2(36),PARTIAL_PRODUCT_2_2(36),PARTIAL_PRODUCT_5_3(36),PARTIAL_PRODUCT_2_3(37));
FA_6_7_8_37_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(37),PARTIAL_PRODUCT_7_2(37),PARTIAL_PRODUCT_8_2(37),PARTIAL_PRODUCT_3_3(37),PARTIAL_PRODUCT_0_3(38));
FA_3_4_5_37_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(37),PARTIAL_PRODUCT_4_2(37),PARTIAL_PRODUCT_5_2(37),PARTIAL_PRODUCT_4_3(37),PARTIAL_PRODUCT_1_3(38));
FA_0_1_2_37_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(37),PARTIAL_PRODUCT_1_2(37),PARTIAL_PRODUCT_2_2(37),PARTIAL_PRODUCT_5_3(37),PARTIAL_PRODUCT_2_3(38));
FA_6_7_8_38_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(38),PARTIAL_PRODUCT_7_2(38),PARTIAL_PRODUCT_8_2(38),PARTIAL_PRODUCT_3_3(38),PARTIAL_PRODUCT_0_3(39));
FA_3_4_5_38_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(38),PARTIAL_PRODUCT_4_2(38),PARTIAL_PRODUCT_5_2(38),PARTIAL_PRODUCT_4_3(38),PARTIAL_PRODUCT_1_3(39));
FA_0_1_2_38_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(38),PARTIAL_PRODUCT_1_2(38),PARTIAL_PRODUCT_2_2(38),PARTIAL_PRODUCT_5_3(38),PARTIAL_PRODUCT_2_3(39));
FA_6_7_8_39_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(39),PARTIAL_PRODUCT_7_2(39),PARTIAL_PRODUCT_8_2(39),PARTIAL_PRODUCT_3_3(39),PARTIAL_PRODUCT_0_3(40));
FA_3_4_5_39_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(39),PARTIAL_PRODUCT_4_2(39),PARTIAL_PRODUCT_5_2(39),PARTIAL_PRODUCT_4_3(39),PARTIAL_PRODUCT_1_3(40));
FA_0_1_2_39_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(39),PARTIAL_PRODUCT_1_2(39),PARTIAL_PRODUCT_2_2(39),PARTIAL_PRODUCT_5_3(39),PARTIAL_PRODUCT_2_3(40));
FA_6_7_8_40_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(40),PARTIAL_PRODUCT_7_2(40),PARTIAL_PRODUCT_8_2(40),PARTIAL_PRODUCT_3_3(40),PARTIAL_PRODUCT_0_3(41));
FA_3_4_5_40_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(40),PARTIAL_PRODUCT_4_2(40),PARTIAL_PRODUCT_5_2(40),PARTIAL_PRODUCT_4_3(40),PARTIAL_PRODUCT_1_3(41));
FA_0_1_2_40_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(40),PARTIAL_PRODUCT_1_2(40),PARTIAL_PRODUCT_2_2(40),PARTIAL_PRODUCT_5_3(40),PARTIAL_PRODUCT_2_3(41));
FA_6_7_8_41_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(41),PARTIAL_PRODUCT_7_2(41),PARTIAL_PRODUCT_8_2(41),PARTIAL_PRODUCT_3_3(41),PARTIAL_PRODUCT_0_3(42));
FA_3_4_5_41_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(41),PARTIAL_PRODUCT_4_2(41),PARTIAL_PRODUCT_5_2(41),PARTIAL_PRODUCT_4_3(41),PARTIAL_PRODUCT_1_3(42));
FA_0_1_2_41_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(41),PARTIAL_PRODUCT_1_2(41),PARTIAL_PRODUCT_2_2(41),PARTIAL_PRODUCT_5_3(41),PARTIAL_PRODUCT_2_3(42));
FA_6_7_8_42_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(42),PARTIAL_PRODUCT_7_2(42),PARTIAL_PRODUCT_8_2(42),PARTIAL_PRODUCT_3_3(42),PARTIAL_PRODUCT_0_3(43));
FA_3_4_5_42_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(42),PARTIAL_PRODUCT_4_2(42),PARTIAL_PRODUCT_5_2(42),PARTIAL_PRODUCT_4_3(42),PARTIAL_PRODUCT_1_3(43));
FA_0_1_2_42_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(42),PARTIAL_PRODUCT_1_2(42),PARTIAL_PRODUCT_2_2(42),PARTIAL_PRODUCT_5_3(42),PARTIAL_PRODUCT_2_3(43));
FA_6_7_8_43_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(43),PARTIAL_PRODUCT_7_2(43),PARTIAL_PRODUCT_8_2(43),PARTIAL_PRODUCT_3_3(43),PARTIAL_PRODUCT_0_3(44));
FA_3_4_5_43_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(43),PARTIAL_PRODUCT_4_2(43),PARTIAL_PRODUCT_5_2(43),PARTIAL_PRODUCT_4_3(43),PARTIAL_PRODUCT_1_3(44));
FA_0_1_2_43_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(43),PARTIAL_PRODUCT_1_2(43),PARTIAL_PRODUCT_2_2(43),PARTIAL_PRODUCT_5_3(43),PARTIAL_PRODUCT_2_3(44));
FA_6_7_8_44_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(44),PARTIAL_PRODUCT_7_2(44),PARTIAL_PRODUCT_8_2(44),PARTIAL_PRODUCT_3_3(44),PARTIAL_PRODUCT_0_3(45));
FA_3_4_5_44_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(44),PARTIAL_PRODUCT_4_2(44),PARTIAL_PRODUCT_5_2(44),PARTIAL_PRODUCT_4_3(44),PARTIAL_PRODUCT_1_3(45));
FA_0_1_2_44_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(44),PARTIAL_PRODUCT_1_2(44),PARTIAL_PRODUCT_2_2(44),PARTIAL_PRODUCT_5_3(44),PARTIAL_PRODUCT_2_3(45));
FA_6_7_8_45_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(45),PARTIAL_PRODUCT_7_2(45),PARTIAL_PRODUCT_8_2(45),PARTIAL_PRODUCT_3_3(45),PARTIAL_PRODUCT_0_3(46));
FA_3_4_5_45_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(45),PARTIAL_PRODUCT_4_2(45),PARTIAL_PRODUCT_5_2(45),PARTIAL_PRODUCT_4_3(45),PARTIAL_PRODUCT_1_3(46));
FA_0_1_2_45_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(45),PARTIAL_PRODUCT_1_2(45),PARTIAL_PRODUCT_2_2(45),PARTIAL_PRODUCT_5_3(45),PARTIAL_PRODUCT_2_3(46));
FA_6_7_8_46_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(46),PARTIAL_PRODUCT_7_2(46),PARTIAL_PRODUCT_8_2(46),PARTIAL_PRODUCT_3_3(46),PARTIAL_PRODUCT_0_3(47));
FA_3_4_5_46_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(46),PARTIAL_PRODUCT_4_2(46),PARTIAL_PRODUCT_5_2(46),PARTIAL_PRODUCT_4_3(46),PARTIAL_PRODUCT_1_3(47));
FA_0_1_2_46_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(46),PARTIAL_PRODUCT_1_2(46),PARTIAL_PRODUCT_2_2(46),PARTIAL_PRODUCT_5_3(46),PARTIAL_PRODUCT_2_3(47));
FA_6_7_8_47_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(47),PARTIAL_PRODUCT_7_2(47),PARTIAL_PRODUCT_8_2(47),PARTIAL_PRODUCT_3_3(47),PARTIAL_PRODUCT_0_3(48));
FA_3_4_5_47_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(47),PARTIAL_PRODUCT_4_2(47),PARTIAL_PRODUCT_5_2(47),PARTIAL_PRODUCT_4_3(47),PARTIAL_PRODUCT_1_3(48));
FA_0_1_2_47_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(47),PARTIAL_PRODUCT_1_2(47),PARTIAL_PRODUCT_2_2(47),PARTIAL_PRODUCT_5_3(47),PARTIAL_PRODUCT_2_3(48));
FA_6_7_8_48_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(48),PARTIAL_PRODUCT_7_2(48),PARTIAL_PRODUCT_8_2(48),PARTIAL_PRODUCT_3_3(48),PARTIAL_PRODUCT_0_3(49));
FA_3_4_5_48_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(48),PARTIAL_PRODUCT_4_2(48),PARTIAL_PRODUCT_5_2(48),PARTIAL_PRODUCT_4_3(48),PARTIAL_PRODUCT_1_3(49));
FA_0_1_2_48_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(48),PARTIAL_PRODUCT_1_2(48),PARTIAL_PRODUCT_2_2(48),PARTIAL_PRODUCT_5_3(48),PARTIAL_PRODUCT_2_3(49));
FA_6_7_8_49_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(49),PARTIAL_PRODUCT_7_2(49),PARTIAL_PRODUCT_8_2(49),PARTIAL_PRODUCT_3_3(49),PARTIAL_PRODUCT_0_3(50));
FA_3_4_5_49_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(49),PARTIAL_PRODUCT_4_2(49),PARTIAL_PRODUCT_5_2(49),PARTIAL_PRODUCT_4_3(49),PARTIAL_PRODUCT_1_3(50));
FA_0_1_2_49_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(49),PARTIAL_PRODUCT_1_2(49),PARTIAL_PRODUCT_2_2(49),PARTIAL_PRODUCT_5_3(49),PARTIAL_PRODUCT_2_3(50));
FA_6_7_8_50_3: FA PORT MAP (PARTIAL_PRODUCT_6_2(50),PARTIAL_PRODUCT_7_2(50),PARTIAL_PRODUCT_8_2(50),PARTIAL_PRODUCT_3_3(50),PARTIAL_PRODUCT_0_3(51));
FA_3_4_5_50_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(50),PARTIAL_PRODUCT_4_2(50),PARTIAL_PRODUCT_5_2(50),PARTIAL_PRODUCT_4_3(50),PARTIAL_PRODUCT_1_3(51));
FA_0_1_2_50_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(50),PARTIAL_PRODUCT_1_2(50),PARTIAL_PRODUCT_2_2(50),PARTIAL_PRODUCT_5_3(50),PARTIAL_PRODUCT_2_3(51));
HA_6_7_51_3: HA PORT MAP (PARTIAL_PRODUCT_6_2(51),PARTIAL_PRODUCT_7_2(51),PARTIAL_PRODUCT_3_3(51),PARTIAL_PRODUCT_0_3(52));
FA_3_4_5_51_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(51),PARTIAL_PRODUCT_4_2(51),PARTIAL_PRODUCT_5_2(51),PARTIAL_PRODUCT_4_3(51),PARTIAL_PRODUCT_1_3(52));
FA_0_1_2_51_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(51),PARTIAL_PRODUCT_1_2(51),PARTIAL_PRODUCT_2_2(51),PARTIAL_PRODUCT_5_3(51),PARTIAL_PRODUCT_2_3(52));
HA_6_7_52_3: HA PORT MAP (PARTIAL_PRODUCT_6_2(52),PARTIAL_PRODUCT_7_2(52),PARTIAL_PRODUCT_3_3(52),PARTIAL_PRODUCT_1_3(53));
FA_3_4_5_52_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(52),PARTIAL_PRODUCT_4_2(52),PARTIAL_PRODUCT_5_2(52),PARTIAL_PRODUCT_4_3(52),PARTIAL_PRODUCT_2_3(53));
FA_0_1_2_52_3: FA PORT MAP (PARTIAL_PRODUCT_0_2(52),PARTIAL_PRODUCT_1_2(52),PARTIAL_PRODUCT_2_2(52),PARTIAL_PRODUCT_5_3(52),PARTIAL_PRODUCT_3_3(53));
FA_4_5_6_53_3: FA PORT MAP (PARTIAL_PRODUCT_4_2(53),PARTIAL_PRODUCT_5_2(53),PARTIAL_PRODUCT_6_2(53),PARTIAL_PRODUCT_4_3(53),PARTIAL_PRODUCT_2_3(54));
FA_1_2_3_53_3: FA PORT MAP (PARTIAL_PRODUCT_1_2(53),PARTIAL_PRODUCT_2_2(53),PARTIAL_PRODUCT_3_2(53),PARTIAL_PRODUCT_5_3(53),PARTIAL_PRODUCT_3_3(54));
HA_5_6_54_3: HA PORT MAP (PARTIAL_PRODUCT_5_2(54),PARTIAL_PRODUCT_6_2(54),PARTIAL_PRODUCT_4_3(54),PARTIAL_PRODUCT_3_3(55));
FA_2_3_4_54_3: FA PORT MAP (PARTIAL_PRODUCT_2_2(54),PARTIAL_PRODUCT_3_2(54),PARTIAL_PRODUCT_4_2(54),PARTIAL_PRODUCT_5_3(54),PARTIAL_PRODUCT_4_3(55));
FA_3_4_5_55_3: FA PORT MAP (PARTIAL_PRODUCT_3_2(55),PARTIAL_PRODUCT_4_2(55),PARTIAL_PRODUCT_5_2(55),PARTIAL_PRODUCT_5_3(55),PARTIAL_PRODUCT_4_3(56));
HA_4_5_56_3: HA PORT MAP (PARTIAL_PRODUCT_4_2(56),PARTIAL_PRODUCT_5_2(56),PARTIAL_PRODUCT_5_3(56),PARTIAL_PRODUCT_5_3(57));


PARTIAL_PRODUCT_0_3( 14 downto 0) <= PARTIAL_PRODUCT_0_2(14 downto 0); 
PARTIAL_PRODUCT_1_3( 13 downto 0) <= PARTIAL_PRODUCT_1_2(13 downto 0); 
PARTIAL_PRODUCT_2_3( 12 downto 0) <= PARTIAL_PRODUCT_2_2(12 downto 0); 
PARTIAL_PRODUCT_3_3( 11 downto 0) <= PARTIAL_PRODUCT_3_2(11 downto 0); 
PARTIAL_PRODUCT_4_3( 10 downto 0) <= PARTIAL_PRODUCT_4_2(10 downto 0); 
PARTIAL_PRODUCT_5_3( 9 downto 0) <= PARTIAL_PRODUCT_5_2(9 downto 0); 
PARTIAL_PRODUCT_1_3( 63 downto 54) <= PARTIAL_PRODUCT_1_2(63 downto 54); 
PARTIAL_PRODUCT_2_3( 63 downto 55) <= PARTIAL_PRODUCT_2_2(63 downto 55); 
PARTIAL_PRODUCT_3_3( 63 downto 56) <= PARTIAL_PRODUCT_3_2(63 downto 56); 
PARTIAL_PRODUCT_4_3( 63 downto 57) <= PARTIAL_PRODUCT_4_2(63 downto 57); 
PARTIAL_PRODUCT_5_3( 63 downto 58) <= PARTIAL_PRODUCT_5_2(63 downto 58); 
PARTIAL_PRODUCT_0_3( 63 downto 53) <= PARTIAL_PRODUCT_0_2(63 downto 53);

HA_3_4_6_4: HA PORT MAP (PARTIAL_PRODUCT_3_3(6),PARTIAL_PRODUCT_4_3(6),PARTIAL_PRODUCT_3_4(6),PARTIAL_PRODUCT_2_4(7));
HA_2_3_7_4: HA PORT MAP (PARTIAL_PRODUCT_2_3(7),PARTIAL_PRODUCT_3_3(7),PARTIAL_PRODUCT_3_4(7),PARTIAL_PRODUCT_1_4(8));
HA_4_5_8_4: HA PORT MAP (PARTIAL_PRODUCT_4_3(8),PARTIAL_PRODUCT_5_3(8),PARTIAL_PRODUCT_2_4(8),PARTIAL_PRODUCT_0_4(9));
FA_1_2_3_8_4: FA PORT MAP (PARTIAL_PRODUCT_1_3(8),PARTIAL_PRODUCT_2_3(8),PARTIAL_PRODUCT_3_3(8),PARTIAL_PRODUCT_3_4(8),PARTIAL_PRODUCT_1_4(9));
HA_3_4_9_4: HA PORT MAP (PARTIAL_PRODUCT_3_3(9),PARTIAL_PRODUCT_4_3(9),PARTIAL_PRODUCT_2_4(9),PARTIAL_PRODUCT_0_4(10));
FA_0_1_2_9_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(9),PARTIAL_PRODUCT_1_3(9),PARTIAL_PRODUCT_2_3(9),PARTIAL_PRODUCT_3_4(9),PARTIAL_PRODUCT_1_4(10));
FA_3_4_5_10_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(10),PARTIAL_PRODUCT_4_3(10),PARTIAL_PRODUCT_5_3(10),PARTIAL_PRODUCT_2_4(10),PARTIAL_PRODUCT_0_4(11));
FA_0_1_2_10_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(10),PARTIAL_PRODUCT_1_3(10),PARTIAL_PRODUCT_2_3(10),PARTIAL_PRODUCT_3_4(10),PARTIAL_PRODUCT_1_4(11));
FA_3_4_5_11_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(11),PARTIAL_PRODUCT_4_3(11),PARTIAL_PRODUCT_5_3(11),PARTIAL_PRODUCT_2_4(11),PARTIAL_PRODUCT_0_4(12));
FA_0_1_2_11_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(11),PARTIAL_PRODUCT_1_3(11),PARTIAL_PRODUCT_2_3(11),PARTIAL_PRODUCT_3_4(11),PARTIAL_PRODUCT_1_4(12));
FA_3_4_5_12_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(12),PARTIAL_PRODUCT_4_3(12),PARTIAL_PRODUCT_5_3(12),PARTIAL_PRODUCT_2_4(12),PARTIAL_PRODUCT_0_4(13));
FA_0_1_2_12_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(12),PARTIAL_PRODUCT_1_3(12),PARTIAL_PRODUCT_2_3(12),PARTIAL_PRODUCT_3_4(12),PARTIAL_PRODUCT_1_4(13));
FA_3_4_5_13_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(13),PARTIAL_PRODUCT_4_3(13),PARTIAL_PRODUCT_5_3(13),PARTIAL_PRODUCT_2_4(13),PARTIAL_PRODUCT_0_4(14));
FA_0_1_2_13_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(13),PARTIAL_PRODUCT_1_3(13),PARTIAL_PRODUCT_2_3(13),PARTIAL_PRODUCT_3_4(13),PARTIAL_PRODUCT_1_4(14));
FA_3_4_5_14_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(14),PARTIAL_PRODUCT_4_3(14),PARTIAL_PRODUCT_5_3(14),PARTIAL_PRODUCT_2_4(14),PARTIAL_PRODUCT_0_4(15));
FA_0_1_2_14_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(14),PARTIAL_PRODUCT_1_3(14),PARTIAL_PRODUCT_2_3(14),PARTIAL_PRODUCT_3_4(14),PARTIAL_PRODUCT_1_4(15));
FA_3_4_5_15_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(15),PARTIAL_PRODUCT_4_3(15),PARTIAL_PRODUCT_5_3(15),PARTIAL_PRODUCT_2_4(15),PARTIAL_PRODUCT_0_4(16));
FA_0_1_2_15_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(15),PARTIAL_PRODUCT_1_3(15),PARTIAL_PRODUCT_2_3(15),PARTIAL_PRODUCT_3_4(15),PARTIAL_PRODUCT_1_4(16));
FA_3_4_5_16_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(16),PARTIAL_PRODUCT_4_3(16),PARTIAL_PRODUCT_5_3(16),PARTIAL_PRODUCT_2_4(16),PARTIAL_PRODUCT_0_4(17));
FA_0_1_2_16_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(16),PARTIAL_PRODUCT_1_3(16),PARTIAL_PRODUCT_2_3(16),PARTIAL_PRODUCT_3_4(16),PARTIAL_PRODUCT_1_4(17));
FA_3_4_5_17_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(17),PARTIAL_PRODUCT_4_3(17),PARTIAL_PRODUCT_5_3(17),PARTIAL_PRODUCT_2_4(17),PARTIAL_PRODUCT_0_4(18));
FA_0_1_2_17_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(17),PARTIAL_PRODUCT_1_3(17),PARTIAL_PRODUCT_2_3(17),PARTIAL_PRODUCT_3_4(17),PARTIAL_PRODUCT_1_4(18));
FA_3_4_5_18_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(18),PARTIAL_PRODUCT_4_3(18),PARTIAL_PRODUCT_5_3(18),PARTIAL_PRODUCT_2_4(18),PARTIAL_PRODUCT_0_4(19));
FA_0_1_2_18_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(18),PARTIAL_PRODUCT_1_3(18),PARTIAL_PRODUCT_2_3(18),PARTIAL_PRODUCT_3_4(18),PARTIAL_PRODUCT_1_4(19));
FA_3_4_5_19_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(19),PARTIAL_PRODUCT_4_3(19),PARTIAL_PRODUCT_5_3(19),PARTIAL_PRODUCT_2_4(19),PARTIAL_PRODUCT_0_4(20));
FA_0_1_2_19_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(19),PARTIAL_PRODUCT_1_3(19),PARTIAL_PRODUCT_2_3(19),PARTIAL_PRODUCT_3_4(19),PARTIAL_PRODUCT_1_4(20));
FA_3_4_5_20_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(20),PARTIAL_PRODUCT_4_3(20),PARTIAL_PRODUCT_5_3(20),PARTIAL_PRODUCT_2_4(20),PARTIAL_PRODUCT_0_4(21));
FA_0_1_2_20_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(20),PARTIAL_PRODUCT_1_3(20),PARTIAL_PRODUCT_2_3(20),PARTIAL_PRODUCT_3_4(20),PARTIAL_PRODUCT_1_4(21));
FA_3_4_5_21_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(21),PARTIAL_PRODUCT_4_3(21),PARTIAL_PRODUCT_5_3(21),PARTIAL_PRODUCT_2_4(21),PARTIAL_PRODUCT_0_4(22));
FA_0_1_2_21_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(21),PARTIAL_PRODUCT_1_3(21),PARTIAL_PRODUCT_2_3(21),PARTIAL_PRODUCT_3_4(21),PARTIAL_PRODUCT_1_4(22));
FA_3_4_5_22_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(22),PARTIAL_PRODUCT_4_3(22),PARTIAL_PRODUCT_5_3(22),PARTIAL_PRODUCT_2_4(22),PARTIAL_PRODUCT_0_4(23));
FA_0_1_2_22_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(22),PARTIAL_PRODUCT_1_3(22),PARTIAL_PRODUCT_2_3(22),PARTIAL_PRODUCT_3_4(22),PARTIAL_PRODUCT_1_4(23));
FA_3_4_5_23_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(23),PARTIAL_PRODUCT_4_3(23),PARTIAL_PRODUCT_5_3(23),PARTIAL_PRODUCT_2_4(23),PARTIAL_PRODUCT_0_4(24));
FA_0_1_2_23_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(23),PARTIAL_PRODUCT_1_3(23),PARTIAL_PRODUCT_2_3(23),PARTIAL_PRODUCT_3_4(23),PARTIAL_PRODUCT_1_4(24));
FA_3_4_5_24_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(24),PARTIAL_PRODUCT_4_3(24),PARTIAL_PRODUCT_5_3(24),PARTIAL_PRODUCT_2_4(24),PARTIAL_PRODUCT_0_4(25));
FA_0_1_2_24_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(24),PARTIAL_PRODUCT_1_3(24),PARTIAL_PRODUCT_2_3(24),PARTIAL_PRODUCT_3_4(24),PARTIAL_PRODUCT_1_4(25));
FA_3_4_5_25_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(25),PARTIAL_PRODUCT_4_3(25),PARTIAL_PRODUCT_5_3(25),PARTIAL_PRODUCT_2_4(25),PARTIAL_PRODUCT_0_4(26));
FA_0_1_2_25_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(25),PARTIAL_PRODUCT_1_3(25),PARTIAL_PRODUCT_2_3(25),PARTIAL_PRODUCT_3_4(25),PARTIAL_PRODUCT_1_4(26));
FA_3_4_5_26_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(26),PARTIAL_PRODUCT_4_3(26),PARTIAL_PRODUCT_5_3(26),PARTIAL_PRODUCT_2_4(26),PARTIAL_PRODUCT_0_4(27));
FA_0_1_2_26_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(26),PARTIAL_PRODUCT_1_3(26),PARTIAL_PRODUCT_2_3(26),PARTIAL_PRODUCT_3_4(26),PARTIAL_PRODUCT_1_4(27));
FA_3_4_5_27_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(27),PARTIAL_PRODUCT_4_3(27),PARTIAL_PRODUCT_5_3(27),PARTIAL_PRODUCT_2_4(27),PARTIAL_PRODUCT_0_4(28));
FA_0_1_2_27_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(27),PARTIAL_PRODUCT_1_3(27),PARTIAL_PRODUCT_2_3(27),PARTIAL_PRODUCT_3_4(27),PARTIAL_PRODUCT_1_4(28));
FA_3_4_5_28_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(28),PARTIAL_PRODUCT_4_3(28),PARTIAL_PRODUCT_5_3(28),PARTIAL_PRODUCT_2_4(28),PARTIAL_PRODUCT_0_4(29));
FA_0_1_2_28_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(28),PARTIAL_PRODUCT_1_3(28),PARTIAL_PRODUCT_2_3(28),PARTIAL_PRODUCT_3_4(28),PARTIAL_PRODUCT_1_4(29));
FA_3_4_5_29_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(29),PARTIAL_PRODUCT_4_3(29),PARTIAL_PRODUCT_5_3(29),PARTIAL_PRODUCT_2_4(29),PARTIAL_PRODUCT_0_4(30));
FA_0_1_2_29_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(29),PARTIAL_PRODUCT_1_3(29),PARTIAL_PRODUCT_2_3(29),PARTIAL_PRODUCT_3_4(29),PARTIAL_PRODUCT_1_4(30));
FA_3_4_5_30_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(30),PARTIAL_PRODUCT_4_3(30),PARTIAL_PRODUCT_5_3(30),PARTIAL_PRODUCT_2_4(30),PARTIAL_PRODUCT_0_4(31));
FA_0_1_2_30_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(30),PARTIAL_PRODUCT_1_3(30),PARTIAL_PRODUCT_2_3(30),PARTIAL_PRODUCT_3_4(30),PARTIAL_PRODUCT_1_4(31));
FA_3_4_5_31_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(31),PARTIAL_PRODUCT_4_3(31),PARTIAL_PRODUCT_5_3(31),PARTIAL_PRODUCT_2_4(31),PARTIAL_PRODUCT_0_4(32));
FA_0_1_2_31_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(31),PARTIAL_PRODUCT_1_3(31),PARTIAL_PRODUCT_2_3(31),PARTIAL_PRODUCT_3_4(31),PARTIAL_PRODUCT_1_4(32));
FA_3_4_5_32_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(32),PARTIAL_PRODUCT_4_3(32),PARTIAL_PRODUCT_5_3(32),PARTIAL_PRODUCT_2_4(32),PARTIAL_PRODUCT_0_4(33));
FA_0_1_2_32_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(32),PARTIAL_PRODUCT_1_3(32),PARTIAL_PRODUCT_2_3(32),PARTIAL_PRODUCT_3_4(32),PARTIAL_PRODUCT_1_4(33));
FA_3_4_5_33_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(33),PARTIAL_PRODUCT_4_3(33),PARTIAL_PRODUCT_5_3(33),PARTIAL_PRODUCT_2_4(33),PARTIAL_PRODUCT_0_4(34));
FA_0_1_2_33_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(33),PARTIAL_PRODUCT_1_3(33),PARTIAL_PRODUCT_2_3(33),PARTIAL_PRODUCT_3_4(33),PARTIAL_PRODUCT_1_4(34));
FA_3_4_5_34_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(34),PARTIAL_PRODUCT_4_3(34),PARTIAL_PRODUCT_5_3(34),PARTIAL_PRODUCT_2_4(34),PARTIAL_PRODUCT_0_4(35));
FA_0_1_2_34_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(34),PARTIAL_PRODUCT_1_3(34),PARTIAL_PRODUCT_2_3(34),PARTIAL_PRODUCT_3_4(34),PARTIAL_PRODUCT_1_4(35));
FA_3_4_5_35_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(35),PARTIAL_PRODUCT_4_3(35),PARTIAL_PRODUCT_5_3(35),PARTIAL_PRODUCT_2_4(35),PARTIAL_PRODUCT_0_4(36));
FA_0_1_2_35_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(35),PARTIAL_PRODUCT_1_3(35),PARTIAL_PRODUCT_2_3(35),PARTIAL_PRODUCT_3_4(35),PARTIAL_PRODUCT_1_4(36));
FA_3_4_5_36_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(36),PARTIAL_PRODUCT_4_3(36),PARTIAL_PRODUCT_5_3(36),PARTIAL_PRODUCT_2_4(36),PARTIAL_PRODUCT_0_4(37));
FA_0_1_2_36_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(36),PARTIAL_PRODUCT_1_3(36),PARTIAL_PRODUCT_2_3(36),PARTIAL_PRODUCT_3_4(36),PARTIAL_PRODUCT_1_4(37));
FA_3_4_5_37_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(37),PARTIAL_PRODUCT_4_3(37),PARTIAL_PRODUCT_5_3(37),PARTIAL_PRODUCT_2_4(37),PARTIAL_PRODUCT_0_4(38));
FA_0_1_2_37_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(37),PARTIAL_PRODUCT_1_3(37),PARTIAL_PRODUCT_2_3(37),PARTIAL_PRODUCT_3_4(37),PARTIAL_PRODUCT_1_4(38));
FA_3_4_5_38_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(38),PARTIAL_PRODUCT_4_3(38),PARTIAL_PRODUCT_5_3(38),PARTIAL_PRODUCT_2_4(38),PARTIAL_PRODUCT_0_4(39));
FA_0_1_2_38_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(38),PARTIAL_PRODUCT_1_3(38),PARTIAL_PRODUCT_2_3(38),PARTIAL_PRODUCT_3_4(38),PARTIAL_PRODUCT_1_4(39));
FA_3_4_5_39_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(39),PARTIAL_PRODUCT_4_3(39),PARTIAL_PRODUCT_5_3(39),PARTIAL_PRODUCT_2_4(39),PARTIAL_PRODUCT_0_4(40));
FA_0_1_2_39_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(39),PARTIAL_PRODUCT_1_3(39),PARTIAL_PRODUCT_2_3(39),PARTIAL_PRODUCT_3_4(39),PARTIAL_PRODUCT_1_4(40));
FA_3_4_5_40_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(40),PARTIAL_PRODUCT_4_3(40),PARTIAL_PRODUCT_5_3(40),PARTIAL_PRODUCT_2_4(40),PARTIAL_PRODUCT_0_4(41));
FA_0_1_2_40_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(40),PARTIAL_PRODUCT_1_3(40),PARTIAL_PRODUCT_2_3(40),PARTIAL_PRODUCT_3_4(40),PARTIAL_PRODUCT_1_4(41));
FA_3_4_5_41_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(41),PARTIAL_PRODUCT_4_3(41),PARTIAL_PRODUCT_5_3(41),PARTIAL_PRODUCT_2_4(41),PARTIAL_PRODUCT_0_4(42));
FA_0_1_2_41_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(41),PARTIAL_PRODUCT_1_3(41),PARTIAL_PRODUCT_2_3(41),PARTIAL_PRODUCT_3_4(41),PARTIAL_PRODUCT_1_4(42));
FA_3_4_5_42_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(42),PARTIAL_PRODUCT_4_3(42),PARTIAL_PRODUCT_5_3(42),PARTIAL_PRODUCT_2_4(42),PARTIAL_PRODUCT_0_4(43));
FA_0_1_2_42_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(42),PARTIAL_PRODUCT_1_3(42),PARTIAL_PRODUCT_2_3(42),PARTIAL_PRODUCT_3_4(42),PARTIAL_PRODUCT_1_4(43));
FA_3_4_5_43_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(43),PARTIAL_PRODUCT_4_3(43),PARTIAL_PRODUCT_5_3(43),PARTIAL_PRODUCT_2_4(43),PARTIAL_PRODUCT_0_4(44));
FA_0_1_2_43_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(43),PARTIAL_PRODUCT_1_3(43),PARTIAL_PRODUCT_2_3(43),PARTIAL_PRODUCT_3_4(43),PARTIAL_PRODUCT_1_4(44));
FA_3_4_5_44_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(44),PARTIAL_PRODUCT_4_3(44),PARTIAL_PRODUCT_5_3(44),PARTIAL_PRODUCT_2_4(44),PARTIAL_PRODUCT_0_4(45));
FA_0_1_2_44_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(44),PARTIAL_PRODUCT_1_3(44),PARTIAL_PRODUCT_2_3(44),PARTIAL_PRODUCT_3_4(44),PARTIAL_PRODUCT_1_4(45));
FA_3_4_5_45_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(45),PARTIAL_PRODUCT_4_3(45),PARTIAL_PRODUCT_5_3(45),PARTIAL_PRODUCT_2_4(45),PARTIAL_PRODUCT_0_4(46));
FA_0_1_2_45_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(45),PARTIAL_PRODUCT_1_3(45),PARTIAL_PRODUCT_2_3(45),PARTIAL_PRODUCT_3_4(45),PARTIAL_PRODUCT_1_4(46));
FA_3_4_5_46_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(46),PARTIAL_PRODUCT_4_3(46),PARTIAL_PRODUCT_5_3(46),PARTIAL_PRODUCT_2_4(46),PARTIAL_PRODUCT_0_4(47));
FA_0_1_2_46_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(46),PARTIAL_PRODUCT_1_3(46),PARTIAL_PRODUCT_2_3(46),PARTIAL_PRODUCT_3_4(46),PARTIAL_PRODUCT_1_4(47));
FA_3_4_5_47_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(47),PARTIAL_PRODUCT_4_3(47),PARTIAL_PRODUCT_5_3(47),PARTIAL_PRODUCT_2_4(47),PARTIAL_PRODUCT_0_4(48));
FA_0_1_2_47_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(47),PARTIAL_PRODUCT_1_3(47),PARTIAL_PRODUCT_2_3(47),PARTIAL_PRODUCT_3_4(47),PARTIAL_PRODUCT_1_4(48));
FA_3_4_5_48_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(48),PARTIAL_PRODUCT_4_3(48),PARTIAL_PRODUCT_5_3(48),PARTIAL_PRODUCT_2_4(48),PARTIAL_PRODUCT_0_4(49));
FA_0_1_2_48_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(48),PARTIAL_PRODUCT_1_3(48),PARTIAL_PRODUCT_2_3(48),PARTIAL_PRODUCT_3_4(48),PARTIAL_PRODUCT_1_4(49));
FA_3_4_5_49_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(49),PARTIAL_PRODUCT_4_3(49),PARTIAL_PRODUCT_5_3(49),PARTIAL_PRODUCT_2_4(49),PARTIAL_PRODUCT_0_4(50));
FA_0_1_2_49_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(49),PARTIAL_PRODUCT_1_3(49),PARTIAL_PRODUCT_2_3(49),PARTIAL_PRODUCT_3_4(49),PARTIAL_PRODUCT_1_4(50));
FA_3_4_5_50_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(50),PARTIAL_PRODUCT_4_3(50),PARTIAL_PRODUCT_5_3(50),PARTIAL_PRODUCT_2_4(50),PARTIAL_PRODUCT_0_4(51));
FA_0_1_2_50_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(50),PARTIAL_PRODUCT_1_3(50),PARTIAL_PRODUCT_2_3(50),PARTIAL_PRODUCT_3_4(50),PARTIAL_PRODUCT_1_4(51));
FA_3_4_5_51_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(51),PARTIAL_PRODUCT_4_3(51),PARTIAL_PRODUCT_5_3(51),PARTIAL_PRODUCT_2_4(51),PARTIAL_PRODUCT_0_4(52));
FA_0_1_2_51_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(51),PARTIAL_PRODUCT_1_3(51),PARTIAL_PRODUCT_2_3(51),PARTIAL_PRODUCT_3_4(51),PARTIAL_PRODUCT_1_4(52));
FA_3_4_5_52_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(52),PARTIAL_PRODUCT_4_3(52),PARTIAL_PRODUCT_5_3(52),PARTIAL_PRODUCT_2_4(52),PARTIAL_PRODUCT_0_4(53));
FA_0_1_2_52_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(52),PARTIAL_PRODUCT_1_3(52),PARTIAL_PRODUCT_2_3(52),PARTIAL_PRODUCT_3_4(52),PARTIAL_PRODUCT_1_4(53));
FA_3_4_5_53_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(53),PARTIAL_PRODUCT_4_3(53),PARTIAL_PRODUCT_5_3(53),PARTIAL_PRODUCT_2_4(53),PARTIAL_PRODUCT_0_4(54));
FA_0_1_2_53_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(53),PARTIAL_PRODUCT_1_3(53),PARTIAL_PRODUCT_2_3(53),PARTIAL_PRODUCT_3_4(53),PARTIAL_PRODUCT_1_4(54));
FA_3_4_5_54_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(54),PARTIAL_PRODUCT_4_3(54),PARTIAL_PRODUCT_5_3(54),PARTIAL_PRODUCT_2_4(54),PARTIAL_PRODUCT_0_4(55));
FA_0_1_2_54_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(54),PARTIAL_PRODUCT_1_3(54),PARTIAL_PRODUCT_2_3(54),PARTIAL_PRODUCT_3_4(54),PARTIAL_PRODUCT_1_4(55));
FA_3_4_5_55_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(55),PARTIAL_PRODUCT_4_3(55),PARTIAL_PRODUCT_5_3(55),PARTIAL_PRODUCT_2_4(55),PARTIAL_PRODUCT_0_4(56));
FA_0_1_2_55_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(55),PARTIAL_PRODUCT_1_3(55),PARTIAL_PRODUCT_2_3(55),PARTIAL_PRODUCT_3_4(55),PARTIAL_PRODUCT_1_4(56));
FA_3_4_5_56_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(56),PARTIAL_PRODUCT_4_3(56),PARTIAL_PRODUCT_5_3(56),PARTIAL_PRODUCT_2_4(56),PARTIAL_PRODUCT_0_4(57));
FA_0_1_2_56_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(56),PARTIAL_PRODUCT_1_3(56),PARTIAL_PRODUCT_2_3(56),PARTIAL_PRODUCT_3_4(56),PARTIAL_PRODUCT_1_4(57));
FA_3_4_5_57_4: FA PORT MAP (PARTIAL_PRODUCT_3_3(57),PARTIAL_PRODUCT_4_3(57),PARTIAL_PRODUCT_5_3(57),PARTIAL_PRODUCT_2_4(57),PARTIAL_PRODUCT_0_4(58));
FA_0_1_2_57_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(57),PARTIAL_PRODUCT_1_3(57),PARTIAL_PRODUCT_2_3(57),PARTIAL_PRODUCT_3_4(57),PARTIAL_PRODUCT_1_4(58));
HA_3_4_58_4: HA PORT MAP (PARTIAL_PRODUCT_3_3(58),PARTIAL_PRODUCT_4_3(58),PARTIAL_PRODUCT_2_4(58),PARTIAL_PRODUCT_1_4(59));
FA_0_1_2_58_4: FA PORT MAP (PARTIAL_PRODUCT_0_3(58),PARTIAL_PRODUCT_1_3(58),PARTIAL_PRODUCT_2_3(58),PARTIAL_PRODUCT_3_4(58),PARTIAL_PRODUCT_2_4(59));
FA_1_2_3_59_4: FA PORT MAP (PARTIAL_PRODUCT_1_3(59),PARTIAL_PRODUCT_2_3(59),PARTIAL_PRODUCT_3_3(59),PARTIAL_PRODUCT_3_4(59),PARTIAL_PRODUCT_2_4(60));
HA_2_3_60_4: HA PORT MAP (PARTIAL_PRODUCT_2_3(60),PARTIAL_PRODUCT_3_3(60),PARTIAL_PRODUCT_3_4(60),PARTIAL_PRODUCT_3_4(61));


PARTIAL_PRODUCT_0_4( 8 downto 0) <= PARTIAL_PRODUCT_0_3(8 downto 0); 
PARTIAL_PRODUCT_1_4( 7 downto 0) <= PARTIAL_PRODUCT_1_3(7 downto 0); 
PARTIAL_PRODUCT_2_4( 6 downto 0) <= PARTIAL_PRODUCT_2_3(6 downto 0); 
PARTIAL_PRODUCT_3_4( 5 downto 0) <= PARTIAL_PRODUCT_3_3(5 downto 0); 
PARTIAL_PRODUCT_0_4( 63 downto 59) <= PARTIAL_PRODUCT_0_3(63 downto 59); 
PARTIAL_PRODUCT_1_4( 63 downto 60) <= PARTIAL_PRODUCT_1_3(63 downto 60); 
PARTIAL_PRODUCT_2_4( 63 downto 61) <= PARTIAL_PRODUCT_2_3(63 downto 61); 
PARTIAL_PRODUCT_3_4( 63 downto 62) <= PARTIAL_PRODUCT_3_3(63 downto 62); 

HA_2_3_4_5: HA PORT MAP (PARTIAL_PRODUCT_2_4(4),PARTIAL_PRODUCT_3_4(4),PARTIAL_PRODUCT_2_5(4),PARTIAL_PRODUCT_1_5(5));
HA_1_2_5_5: HA PORT MAP (PARTIAL_PRODUCT_1_4(5),PARTIAL_PRODUCT_2_4(5),PARTIAL_PRODUCT_2_5(5),PARTIAL_PRODUCT_1_5(6));
FA_1_2_3_6_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(6),PARTIAL_PRODUCT_2_4(6),PARTIAL_PRODUCT_3_4(6),PARTIAL_PRODUCT_2_5(6),PARTIAL_PRODUCT_1_5(7));
FA_1_2_3_7_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(7),PARTIAL_PRODUCT_2_4(7),PARTIAL_PRODUCT_3_4(7),PARTIAL_PRODUCT_2_5(7),PARTIAL_PRODUCT_1_5(8));
FA_1_2_3_8_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(8),PARTIAL_PRODUCT_2_4(8),PARTIAL_PRODUCT_3_4(8),PARTIAL_PRODUCT_2_5(8),PARTIAL_PRODUCT_1_5(9));
FA_1_2_3_9_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(9),PARTIAL_PRODUCT_2_4(9),PARTIAL_PRODUCT_3_4(9),PARTIAL_PRODUCT_2_5(9),PARTIAL_PRODUCT_1_5(10));
FA_1_2_3_10_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(10),PARTIAL_PRODUCT_2_4(10),PARTIAL_PRODUCT_3_4(10),PARTIAL_PRODUCT_2_5(10),PARTIAL_PRODUCT_1_5(11));
FA_1_2_3_11_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(11),PARTIAL_PRODUCT_2_4(11),PARTIAL_PRODUCT_3_4(11),PARTIAL_PRODUCT_2_5(11),PARTIAL_PRODUCT_1_5(12));
FA_1_2_3_12_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(12),PARTIAL_PRODUCT_2_4(12),PARTIAL_PRODUCT_3_4(12),PARTIAL_PRODUCT_2_5(12),PARTIAL_PRODUCT_1_5(13));
FA_1_2_3_13_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(13),PARTIAL_PRODUCT_2_4(13),PARTIAL_PRODUCT_3_4(13),PARTIAL_PRODUCT_2_5(13),PARTIAL_PRODUCT_1_5(14));
FA_1_2_3_14_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(14),PARTIAL_PRODUCT_2_4(14),PARTIAL_PRODUCT_3_4(14),PARTIAL_PRODUCT_2_5(14),PARTIAL_PRODUCT_1_5(15));
FA_1_2_3_15_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(15),PARTIAL_PRODUCT_2_4(15),PARTIAL_PRODUCT_3_4(15),PARTIAL_PRODUCT_2_5(15),PARTIAL_PRODUCT_1_5(16));
FA_1_2_3_16_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(16),PARTIAL_PRODUCT_2_4(16),PARTIAL_PRODUCT_3_4(16),PARTIAL_PRODUCT_2_5(16),PARTIAL_PRODUCT_1_5(17));
FA_1_2_3_17_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(17),PARTIAL_PRODUCT_2_4(17),PARTIAL_PRODUCT_3_4(17),PARTIAL_PRODUCT_2_5(17),PARTIAL_PRODUCT_1_5(18));
FA_1_2_3_18_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(18),PARTIAL_PRODUCT_2_4(18),PARTIAL_PRODUCT_3_4(18),PARTIAL_PRODUCT_2_5(18),PARTIAL_PRODUCT_1_5(19));
FA_1_2_3_19_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(19),PARTIAL_PRODUCT_2_4(19),PARTIAL_PRODUCT_3_4(19),PARTIAL_PRODUCT_2_5(19),PARTIAL_PRODUCT_1_5(20));
FA_1_2_3_20_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(20),PARTIAL_PRODUCT_2_4(20),PARTIAL_PRODUCT_3_4(20),PARTIAL_PRODUCT_2_5(20),PARTIAL_PRODUCT_1_5(21));
FA_1_2_3_21_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(21),PARTIAL_PRODUCT_2_4(21),PARTIAL_PRODUCT_3_4(21),PARTIAL_PRODUCT_2_5(21),PARTIAL_PRODUCT_1_5(22));
FA_1_2_3_22_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(22),PARTIAL_PRODUCT_2_4(22),PARTIAL_PRODUCT_3_4(22),PARTIAL_PRODUCT_2_5(22),PARTIAL_PRODUCT_1_5(23));
FA_1_2_3_23_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(23),PARTIAL_PRODUCT_2_4(23),PARTIAL_PRODUCT_3_4(23),PARTIAL_PRODUCT_2_5(23),PARTIAL_PRODUCT_1_5(24));
FA_1_2_3_24_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(24),PARTIAL_PRODUCT_2_4(24),PARTIAL_PRODUCT_3_4(24),PARTIAL_PRODUCT_2_5(24),PARTIAL_PRODUCT_1_5(25));
FA_1_2_3_25_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(25),PARTIAL_PRODUCT_2_4(25),PARTIAL_PRODUCT_3_4(25),PARTIAL_PRODUCT_2_5(25),PARTIAL_PRODUCT_1_5(26));
FA_1_2_3_26_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(26),PARTIAL_PRODUCT_2_4(26),PARTIAL_PRODUCT_3_4(26),PARTIAL_PRODUCT_2_5(26),PARTIAL_PRODUCT_1_5(27));
FA_1_2_3_27_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(27),PARTIAL_PRODUCT_2_4(27),PARTIAL_PRODUCT_3_4(27),PARTIAL_PRODUCT_2_5(27),PARTIAL_PRODUCT_1_5(28));
FA_1_2_3_28_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(28),PARTIAL_PRODUCT_2_4(28),PARTIAL_PRODUCT_3_4(28),PARTIAL_PRODUCT_2_5(28),PARTIAL_PRODUCT_1_5(29));
FA_1_2_3_29_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(29),PARTIAL_PRODUCT_2_4(29),PARTIAL_PRODUCT_3_4(29),PARTIAL_PRODUCT_2_5(29),PARTIAL_PRODUCT_1_5(30));
FA_1_2_3_30_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(30),PARTIAL_PRODUCT_2_4(30),PARTIAL_PRODUCT_3_4(30),PARTIAL_PRODUCT_2_5(30),PARTIAL_PRODUCT_1_5(31));
FA_1_2_3_31_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(31),PARTIAL_PRODUCT_2_4(31),PARTIAL_PRODUCT_3_4(31),PARTIAL_PRODUCT_2_5(31),PARTIAL_PRODUCT_1_5(32));
FA_1_2_3_32_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(32),PARTIAL_PRODUCT_2_4(32),PARTIAL_PRODUCT_3_4(32),PARTIAL_PRODUCT_2_5(32),PARTIAL_PRODUCT_1_5(33));
FA_1_2_3_33_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(33),PARTIAL_PRODUCT_2_4(33),PARTIAL_PRODUCT_3_4(33),PARTIAL_PRODUCT_2_5(33),PARTIAL_PRODUCT_1_5(34));
FA_1_2_3_34_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(34),PARTIAL_PRODUCT_2_4(34),PARTIAL_PRODUCT_3_4(34),PARTIAL_PRODUCT_2_5(34),PARTIAL_PRODUCT_1_5(35));
FA_1_2_3_35_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(35),PARTIAL_PRODUCT_2_4(35),PARTIAL_PRODUCT_3_4(35),PARTIAL_PRODUCT_2_5(35),PARTIAL_PRODUCT_1_5(36));
FA_1_2_3_36_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(36),PARTIAL_PRODUCT_2_4(36),PARTIAL_PRODUCT_3_4(36),PARTIAL_PRODUCT_2_5(36),PARTIAL_PRODUCT_1_5(37));
FA_1_2_3_37_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(37),PARTIAL_PRODUCT_2_4(37),PARTIAL_PRODUCT_3_4(37),PARTIAL_PRODUCT_2_5(37),PARTIAL_PRODUCT_1_5(38));
FA_1_2_3_38_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(38),PARTIAL_PRODUCT_2_4(38),PARTIAL_PRODUCT_3_4(38),PARTIAL_PRODUCT_2_5(38),PARTIAL_PRODUCT_1_5(39));
FA_1_2_3_39_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(39),PARTIAL_PRODUCT_2_4(39),PARTIAL_PRODUCT_3_4(39),PARTIAL_PRODUCT_2_5(39),PARTIAL_PRODUCT_1_5(40));
FA_1_2_3_40_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(40),PARTIAL_PRODUCT_2_4(40),PARTIAL_PRODUCT_3_4(40),PARTIAL_PRODUCT_2_5(40),PARTIAL_PRODUCT_1_5(41));
FA_1_2_3_41_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(41),PARTIAL_PRODUCT_2_4(41),PARTIAL_PRODUCT_3_4(41),PARTIAL_PRODUCT_2_5(41),PARTIAL_PRODUCT_1_5(42));
FA_1_2_3_42_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(42),PARTIAL_PRODUCT_2_4(42),PARTIAL_PRODUCT_3_4(42),PARTIAL_PRODUCT_2_5(42),PARTIAL_PRODUCT_1_5(43));
FA_1_2_3_43_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(43),PARTIAL_PRODUCT_2_4(43),PARTIAL_PRODUCT_3_4(43),PARTIAL_PRODUCT_2_5(43),PARTIAL_PRODUCT_1_5(44));
FA_1_2_3_44_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(44),PARTIAL_PRODUCT_2_4(44),PARTIAL_PRODUCT_3_4(44),PARTIAL_PRODUCT_2_5(44),PARTIAL_PRODUCT_1_5(45));
FA_1_2_3_45_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(45),PARTIAL_PRODUCT_2_4(45),PARTIAL_PRODUCT_3_4(45),PARTIAL_PRODUCT_2_5(45),PARTIAL_PRODUCT_1_5(46));
FA_1_2_3_46_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(46),PARTIAL_PRODUCT_2_4(46),PARTIAL_PRODUCT_3_4(46),PARTIAL_PRODUCT_2_5(46),PARTIAL_PRODUCT_1_5(47));
FA_1_2_3_47_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(47),PARTIAL_PRODUCT_2_4(47),PARTIAL_PRODUCT_3_4(47),PARTIAL_PRODUCT_2_5(47),PARTIAL_PRODUCT_1_5(48));
FA_1_2_3_48_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(48),PARTIAL_PRODUCT_2_4(48),PARTIAL_PRODUCT_3_4(48),PARTIAL_PRODUCT_2_5(48),PARTIAL_PRODUCT_1_5(49));
FA_1_2_3_49_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(49),PARTIAL_PRODUCT_2_4(49),PARTIAL_PRODUCT_3_4(49),PARTIAL_PRODUCT_2_5(49),PARTIAL_PRODUCT_1_5(50));
FA_1_2_3_50_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(50),PARTIAL_PRODUCT_2_4(50),PARTIAL_PRODUCT_3_4(50),PARTIAL_PRODUCT_2_5(50),PARTIAL_PRODUCT_1_5(51));
FA_1_2_3_51_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(51),PARTIAL_PRODUCT_2_4(51),PARTIAL_PRODUCT_3_4(51),PARTIAL_PRODUCT_2_5(51),PARTIAL_PRODUCT_1_5(52));
FA_1_2_3_52_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(52),PARTIAL_PRODUCT_2_4(52),PARTIAL_PRODUCT_3_4(52),PARTIAL_PRODUCT_2_5(52),PARTIAL_PRODUCT_1_5(53));
FA_1_2_3_53_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(53),PARTIAL_PRODUCT_2_4(53),PARTIAL_PRODUCT_3_4(53),PARTIAL_PRODUCT_2_5(53),PARTIAL_PRODUCT_1_5(54));
FA_1_2_3_54_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(54),PARTIAL_PRODUCT_2_4(54),PARTIAL_PRODUCT_3_4(54),PARTIAL_PRODUCT_2_5(54),PARTIAL_PRODUCT_1_5(55));
FA_1_2_3_55_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(55),PARTIAL_PRODUCT_2_4(55),PARTIAL_PRODUCT_3_4(55),PARTIAL_PRODUCT_2_5(55),PARTIAL_PRODUCT_1_5(56));
FA_1_2_3_56_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(56),PARTIAL_PRODUCT_2_4(56),PARTIAL_PRODUCT_3_4(56),PARTIAL_PRODUCT_2_5(56),PARTIAL_PRODUCT_1_5(57));
FA_1_2_3_57_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(57),PARTIAL_PRODUCT_2_4(57),PARTIAL_PRODUCT_3_4(57),PARTIAL_PRODUCT_2_5(57),PARTIAL_PRODUCT_1_5(58));
FA_1_2_3_58_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(58),PARTIAL_PRODUCT_2_4(58),PARTIAL_PRODUCT_3_4(58),PARTIAL_PRODUCT_2_5(58),PARTIAL_PRODUCT_1_5(59));
FA_1_2_3_59_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(59),PARTIAL_PRODUCT_2_4(59),PARTIAL_PRODUCT_3_4(59),PARTIAL_PRODUCT_2_5(59),PARTIAL_PRODUCT_1_5(60));
FA_1_2_3_60_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(60),PARTIAL_PRODUCT_2_4(60),PARTIAL_PRODUCT_3_4(60),PARTIAL_PRODUCT_2_5(60),PARTIAL_PRODUCT_1_5(61));
FA_1_2_3_61_5: FA PORT MAP (PARTIAL_PRODUCT_1_4(61),PARTIAL_PRODUCT_2_4(61),PARTIAL_PRODUCT_3_4(61),PARTIAL_PRODUCT_2_5(61),PARTIAL_PRODUCT_1_5(62));
HA_1_2_62_5: HA PORT MAP (PARTIAL_PRODUCT_1_4(62),PARTIAL_PRODUCT_2_4(62),PARTIAL_PRODUCT_2_5(62),PARTIAL_PRODUCT_2_5(63));



PARTIAL_PRODUCT_0_5( 63 downto 0) <= PARTIAL_PRODUCT_0_4(63 downto 0); 
PARTIAL_PRODUCT_1_5( 4 downto 0) <= PARTIAL_PRODUCT_1_4(4 downto 0); 
PARTIAL_PRODUCT_2_5( 3 downto 0) <= PARTIAL_PRODUCT_2_4(3 downto 0); 
PARTIAL_PRODUCT_1_5( 63 downto 63) <= PARTIAL_PRODUCT_1_4(63 downto 63); 

HA_1_2_2_6: HA PORT MAP (PARTIAL_PRODUCT_1_5(2),PARTIAL_PRODUCT_2_5(2),PARTIAL_PRODUCT_1_6(2),PARTIAL_PRODUCT_0_6(3));
HA_0_1_3_6: HA PORT MAP (PARTIAL_PRODUCT_0_5(3),PARTIAL_PRODUCT_1_5(3),PARTIAL_PRODUCT_1_6(3),PARTIAL_PRODUCT_0_6(4));
FA_0_1_2_4_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(4),PARTIAL_PRODUCT_1_5(4),PARTIAL_PRODUCT_2_5(4),PARTIAL_PRODUCT_1_6(4),PARTIAL_PRODUCT_0_6(5));
FA_0_1_2_5_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(5),PARTIAL_PRODUCT_1_5(5),PARTIAL_PRODUCT_2_5(5),PARTIAL_PRODUCT_1_6(5),PARTIAL_PRODUCT_0_6(6));
FA_0_1_2_6_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(6),PARTIAL_PRODUCT_1_5(6),PARTIAL_PRODUCT_2_5(6),PARTIAL_PRODUCT_1_6(6),PARTIAL_PRODUCT_0_6(7));
FA_0_1_2_7_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(7),PARTIAL_PRODUCT_1_5(7),PARTIAL_PRODUCT_2_5(7),PARTIAL_PRODUCT_1_6(7),PARTIAL_PRODUCT_0_6(8));
FA_0_1_2_8_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(8),PARTIAL_PRODUCT_1_5(8),PARTIAL_PRODUCT_2_5(8),PARTIAL_PRODUCT_1_6(8),PARTIAL_PRODUCT_0_6(9));
FA_0_1_2_9_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(9),PARTIAL_PRODUCT_1_5(9),PARTIAL_PRODUCT_2_5(9),PARTIAL_PRODUCT_1_6(9),PARTIAL_PRODUCT_0_6(10));
FA_0_1_2_10_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(10),PARTIAL_PRODUCT_1_5(10),PARTIAL_PRODUCT_2_5(10),PARTIAL_PRODUCT_1_6(10),PARTIAL_PRODUCT_0_6(11));
FA_0_1_2_11_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(11),PARTIAL_PRODUCT_1_5(11),PARTIAL_PRODUCT_2_5(11),PARTIAL_PRODUCT_1_6(11),PARTIAL_PRODUCT_0_6(12));
FA_0_1_2_12_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(12),PARTIAL_PRODUCT_1_5(12),PARTIAL_PRODUCT_2_5(12),PARTIAL_PRODUCT_1_6(12),PARTIAL_PRODUCT_0_6(13));
FA_0_1_2_13_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(13),PARTIAL_PRODUCT_1_5(13),PARTIAL_PRODUCT_2_5(13),PARTIAL_PRODUCT_1_6(13),PARTIAL_PRODUCT_0_6(14));
FA_0_1_2_14_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(14),PARTIAL_PRODUCT_1_5(14),PARTIAL_PRODUCT_2_5(14),PARTIAL_PRODUCT_1_6(14),PARTIAL_PRODUCT_0_6(15));
FA_0_1_2_15_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(15),PARTIAL_PRODUCT_1_5(15),PARTIAL_PRODUCT_2_5(15),PARTIAL_PRODUCT_1_6(15),PARTIAL_PRODUCT_0_6(16));
FA_0_1_2_16_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(16),PARTIAL_PRODUCT_1_5(16),PARTIAL_PRODUCT_2_5(16),PARTIAL_PRODUCT_1_6(16),PARTIAL_PRODUCT_0_6(17));
FA_0_1_2_17_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(17),PARTIAL_PRODUCT_1_5(17),PARTIAL_PRODUCT_2_5(17),PARTIAL_PRODUCT_1_6(17),PARTIAL_PRODUCT_0_6(18));
FA_0_1_2_18_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(18),PARTIAL_PRODUCT_1_5(18),PARTIAL_PRODUCT_2_5(18),PARTIAL_PRODUCT_1_6(18),PARTIAL_PRODUCT_0_6(19));
FA_0_1_2_19_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(19),PARTIAL_PRODUCT_1_5(19),PARTIAL_PRODUCT_2_5(19),PARTIAL_PRODUCT_1_6(19),PARTIAL_PRODUCT_0_6(20));
FA_0_1_2_20_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(20),PARTIAL_PRODUCT_1_5(20),PARTIAL_PRODUCT_2_5(20),PARTIAL_PRODUCT_1_6(20),PARTIAL_PRODUCT_0_6(21));
FA_0_1_2_21_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(21),PARTIAL_PRODUCT_1_5(21),PARTIAL_PRODUCT_2_5(21),PARTIAL_PRODUCT_1_6(21),PARTIAL_PRODUCT_0_6(22));
FA_0_1_2_22_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(22),PARTIAL_PRODUCT_1_5(22),PARTIAL_PRODUCT_2_5(22),PARTIAL_PRODUCT_1_6(22),PARTIAL_PRODUCT_0_6(23));
FA_0_1_2_23_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(23),PARTIAL_PRODUCT_1_5(23),PARTIAL_PRODUCT_2_5(23),PARTIAL_PRODUCT_1_6(23),PARTIAL_PRODUCT_0_6(24));
FA_0_1_2_24_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(24),PARTIAL_PRODUCT_1_5(24),PARTIAL_PRODUCT_2_5(24),PARTIAL_PRODUCT_1_6(24),PARTIAL_PRODUCT_0_6(25));
FA_0_1_2_25_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(25),PARTIAL_PRODUCT_1_5(25),PARTIAL_PRODUCT_2_5(25),PARTIAL_PRODUCT_1_6(25),PARTIAL_PRODUCT_0_6(26));
FA_0_1_2_26_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(26),PARTIAL_PRODUCT_1_5(26),PARTIAL_PRODUCT_2_5(26),PARTIAL_PRODUCT_1_6(26),PARTIAL_PRODUCT_0_6(27));
FA_0_1_2_27_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(27),PARTIAL_PRODUCT_1_5(27),PARTIAL_PRODUCT_2_5(27),PARTIAL_PRODUCT_1_6(27),PARTIAL_PRODUCT_0_6(28));
FA_0_1_2_28_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(28),PARTIAL_PRODUCT_1_5(28),PARTIAL_PRODUCT_2_5(28),PARTIAL_PRODUCT_1_6(28),PARTIAL_PRODUCT_0_6(29));
FA_0_1_2_29_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(29),PARTIAL_PRODUCT_1_5(29),PARTIAL_PRODUCT_2_5(29),PARTIAL_PRODUCT_1_6(29),PARTIAL_PRODUCT_0_6(30));
FA_0_1_2_30_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(30),PARTIAL_PRODUCT_1_5(30),PARTIAL_PRODUCT_2_5(30),PARTIAL_PRODUCT_1_6(30),PARTIAL_PRODUCT_0_6(31));
FA_0_1_2_31_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(31),PARTIAL_PRODUCT_1_5(31),PARTIAL_PRODUCT_2_5(31),PARTIAL_PRODUCT_1_6(31),PARTIAL_PRODUCT_0_6(32));
FA_0_1_2_32_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(32),PARTIAL_PRODUCT_1_5(32),PARTIAL_PRODUCT_2_5(32),PARTIAL_PRODUCT_1_6(32),PARTIAL_PRODUCT_0_6(33));
FA_0_1_2_33_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(33),PARTIAL_PRODUCT_1_5(33),PARTIAL_PRODUCT_2_5(33),PARTIAL_PRODUCT_1_6(33),PARTIAL_PRODUCT_0_6(34));
FA_0_1_2_34_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(34),PARTIAL_PRODUCT_1_5(34),PARTIAL_PRODUCT_2_5(34),PARTIAL_PRODUCT_1_6(34),PARTIAL_PRODUCT_0_6(35));
FA_0_1_2_35_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(35),PARTIAL_PRODUCT_1_5(35),PARTIAL_PRODUCT_2_5(35),PARTIAL_PRODUCT_1_6(35),PARTIAL_PRODUCT_0_6(36));
FA_0_1_2_36_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(36),PARTIAL_PRODUCT_1_5(36),PARTIAL_PRODUCT_2_5(36),PARTIAL_PRODUCT_1_6(36),PARTIAL_PRODUCT_0_6(37));
FA_0_1_2_37_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(37),PARTIAL_PRODUCT_1_5(37),PARTIAL_PRODUCT_2_5(37),PARTIAL_PRODUCT_1_6(37),PARTIAL_PRODUCT_0_6(38));
FA_0_1_2_38_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(38),PARTIAL_PRODUCT_1_5(38),PARTIAL_PRODUCT_2_5(38),PARTIAL_PRODUCT_1_6(38),PARTIAL_PRODUCT_0_6(39));
FA_0_1_2_39_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(39),PARTIAL_PRODUCT_1_5(39),PARTIAL_PRODUCT_2_5(39),PARTIAL_PRODUCT_1_6(39),PARTIAL_PRODUCT_0_6(40));
FA_0_1_2_40_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(40),PARTIAL_PRODUCT_1_5(40),PARTIAL_PRODUCT_2_5(40),PARTIAL_PRODUCT_1_6(40),PARTIAL_PRODUCT_0_6(41));
FA_0_1_2_41_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(41),PARTIAL_PRODUCT_1_5(41),PARTIAL_PRODUCT_2_5(41),PARTIAL_PRODUCT_1_6(41),PARTIAL_PRODUCT_0_6(42));
FA_0_1_2_42_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(42),PARTIAL_PRODUCT_1_5(42),PARTIAL_PRODUCT_2_5(42),PARTIAL_PRODUCT_1_6(42),PARTIAL_PRODUCT_0_6(43));
FA_0_1_2_43_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(43),PARTIAL_PRODUCT_1_5(43),PARTIAL_PRODUCT_2_5(43),PARTIAL_PRODUCT_1_6(43),PARTIAL_PRODUCT_0_6(44));
FA_0_1_2_44_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(44),PARTIAL_PRODUCT_1_5(44),PARTIAL_PRODUCT_2_5(44),PARTIAL_PRODUCT_1_6(44),PARTIAL_PRODUCT_0_6(45));
FA_0_1_2_45_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(45),PARTIAL_PRODUCT_1_5(45),PARTIAL_PRODUCT_2_5(45),PARTIAL_PRODUCT_1_6(45),PARTIAL_PRODUCT_0_6(46));
FA_0_1_2_46_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(46),PARTIAL_PRODUCT_1_5(46),PARTIAL_PRODUCT_2_5(46),PARTIAL_PRODUCT_1_6(46),PARTIAL_PRODUCT_0_6(47));
FA_0_1_2_47_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(47),PARTIAL_PRODUCT_1_5(47),PARTIAL_PRODUCT_2_5(47),PARTIAL_PRODUCT_1_6(47),PARTIAL_PRODUCT_0_6(48));
FA_0_1_2_48_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(48),PARTIAL_PRODUCT_1_5(48),PARTIAL_PRODUCT_2_5(48),PARTIAL_PRODUCT_1_6(48),PARTIAL_PRODUCT_0_6(49));
FA_0_1_2_49_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(49),PARTIAL_PRODUCT_1_5(49),PARTIAL_PRODUCT_2_5(49),PARTIAL_PRODUCT_1_6(49),PARTIAL_PRODUCT_0_6(50));
FA_0_1_2_50_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(50),PARTIAL_PRODUCT_1_5(50),PARTIAL_PRODUCT_2_5(50),PARTIAL_PRODUCT_1_6(50),PARTIAL_PRODUCT_0_6(51));
FA_0_1_2_51_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(51),PARTIAL_PRODUCT_1_5(51),PARTIAL_PRODUCT_2_5(51),PARTIAL_PRODUCT_1_6(51),PARTIAL_PRODUCT_0_6(52));
FA_0_1_2_52_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(52),PARTIAL_PRODUCT_1_5(52),PARTIAL_PRODUCT_2_5(52),PARTIAL_PRODUCT_1_6(52),PARTIAL_PRODUCT_0_6(53));
FA_0_1_2_53_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(53),PARTIAL_PRODUCT_1_5(53),PARTIAL_PRODUCT_2_5(53),PARTIAL_PRODUCT_1_6(53),PARTIAL_PRODUCT_0_6(54));
FA_0_1_2_54_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(54),PARTIAL_PRODUCT_1_5(54),PARTIAL_PRODUCT_2_5(54),PARTIAL_PRODUCT_1_6(54),PARTIAL_PRODUCT_0_6(55));
FA_0_1_2_55_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(55),PARTIAL_PRODUCT_1_5(55),PARTIAL_PRODUCT_2_5(55),PARTIAL_PRODUCT_1_6(55),PARTIAL_PRODUCT_0_6(56));
FA_0_1_2_56_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(56),PARTIAL_PRODUCT_1_5(56),PARTIAL_PRODUCT_2_5(56),PARTIAL_PRODUCT_1_6(56),PARTIAL_PRODUCT_0_6(57));
FA_0_1_2_57_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(57),PARTIAL_PRODUCT_1_5(57),PARTIAL_PRODUCT_2_5(57),PARTIAL_PRODUCT_1_6(57),PARTIAL_PRODUCT_0_6(58));
FA_0_1_2_58_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(58),PARTIAL_PRODUCT_1_5(58),PARTIAL_PRODUCT_2_5(58),PARTIAL_PRODUCT_1_6(58),PARTIAL_PRODUCT_0_6(59));
FA_0_1_2_59_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(59),PARTIAL_PRODUCT_1_5(59),PARTIAL_PRODUCT_2_5(59),PARTIAL_PRODUCT_1_6(59),PARTIAL_PRODUCT_0_6(60));
FA_0_1_2_60_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(60),PARTIAL_PRODUCT_1_5(60),PARTIAL_PRODUCT_2_5(60),PARTIAL_PRODUCT_1_6(60),PARTIAL_PRODUCT_0_6(61));
FA_0_1_2_61_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(61),PARTIAL_PRODUCT_1_5(61),PARTIAL_PRODUCT_2_5(61),PARTIAL_PRODUCT_1_6(61),PARTIAL_PRODUCT_0_6(62));
FA_0_1_2_62_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(62),PARTIAL_PRODUCT_1_5(62),PARTIAL_PRODUCT_2_5(62),PARTIAL_PRODUCT_1_6(62),PARTIAL_PRODUCT_0_6(63));
FA_0_1_2_63_6: FA PORT MAP (PARTIAL_PRODUCT_0_5(63),PARTIAL_PRODUCT_1_5(63),PARTIAL_PRODUCT_2_5(63),PARTIAL_PRODUCT_1_6(63),CARRY_6);



PARTIAL_PRODUCT_0_6( 2 downto 0) <= PARTIAL_PRODUCT_0_5(2 downto 0); 
PARTIAL_PRODUCT_1_6( 1 downto 0) <= PARTIAL_PRODUCT_1_5(1 downto 0); 
--PARTIAL_PRODUCT_1_6( 63 downto 0) <= PARTIAL_PRODUCT_1_5(63 downto 0); 

HA_0_1_0_7: HA PORT MAP (PARTIAL_PRODUCT_0_6(0),PARTIAL_PRODUCT_1_6(0),PARTIAL_PRODUCT_0_7(0),CARRY_OUT_7(0));
HA_C_0_1_7: HA PORT MAP (CARRY_OUT_7(0),PARTIAL_PRODUCT_0_6(1),PARTIAL_PRODUCT_0_7(1),CARRY_OUT_7(1));
FA_C_0_1_2_7: FA PORT MAP (CARRY_OUT_7(1),PARTIAL_PRODUCT_0_6(2),PARTIAL_PRODUCT_1_6(2),PARTIAL_PRODUCT_0_7(2),CARRY_OUT_7(2));
FA_C_0_1_3_7: FA PORT MAP (CARRY_OUT_7(2),PARTIAL_PRODUCT_0_6(3),PARTIAL_PRODUCT_1_6(3),PARTIAL_PRODUCT_0_7(3),CARRY_OUT_7(3));
FA_C_0_1_4_7: FA PORT MAP (CARRY_OUT_7(3),PARTIAL_PRODUCT_0_6(4),PARTIAL_PRODUCT_1_6(4),PARTIAL_PRODUCT_0_7(4),CARRY_OUT_7(4));
FA_C_0_1_5_7: FA PORT MAP (CARRY_OUT_7(4),PARTIAL_PRODUCT_0_6(5),PARTIAL_PRODUCT_1_6(5),PARTIAL_PRODUCT_0_7(5),CARRY_OUT_7(5));
FA_C_0_1_6_7: FA PORT MAP (CARRY_OUT_7(5),PARTIAL_PRODUCT_0_6(6),PARTIAL_PRODUCT_1_6(6),PARTIAL_PRODUCT_0_7(6),CARRY_OUT_7(6));
FA_C_0_1_7_7: FA PORT MAP (CARRY_OUT_7(6),PARTIAL_PRODUCT_0_6(7),PARTIAL_PRODUCT_1_6(7),PARTIAL_PRODUCT_0_7(7),CARRY_OUT_7(7));
FA_C_0_1_8_7: FA PORT MAP (CARRY_OUT_7(7),PARTIAL_PRODUCT_0_6(8),PARTIAL_PRODUCT_1_6(8),PARTIAL_PRODUCT_0_7(8),CARRY_OUT_7(8));
FA_C_0_1_9_7: FA PORT MAP (CARRY_OUT_7(8),PARTIAL_PRODUCT_0_6(9),PARTIAL_PRODUCT_1_6(9),PARTIAL_PRODUCT_0_7(9),CARRY_OUT_7(9));
FA_C_0_1_10_7: FA PORT MAP (CARRY_OUT_7(9),PARTIAL_PRODUCT_0_6(10),PARTIAL_PRODUCT_1_6(10),PARTIAL_PRODUCT_0_7(10),CARRY_OUT_7(10));
FA_C_0_1_11_7: FA PORT MAP (CARRY_OUT_7(10),PARTIAL_PRODUCT_0_6(11),PARTIAL_PRODUCT_1_6(11),PARTIAL_PRODUCT_0_7(11),CARRY_OUT_7(11));
FA_C_0_1_12_7: FA PORT MAP (CARRY_OUT_7(11),PARTIAL_PRODUCT_0_6(12),PARTIAL_PRODUCT_1_6(12),PARTIAL_PRODUCT_0_7(12),CARRY_OUT_7(12));
FA_C_0_1_13_7: FA PORT MAP (CARRY_OUT_7(12),PARTIAL_PRODUCT_0_6(13),PARTIAL_PRODUCT_1_6(13),PARTIAL_PRODUCT_0_7(13),CARRY_OUT_7(13));
FA_C_0_1_14_7: FA PORT MAP (CARRY_OUT_7(13),PARTIAL_PRODUCT_0_6(14),PARTIAL_PRODUCT_1_6(14),PARTIAL_PRODUCT_0_7(14),CARRY_OUT_7(14));
FA_C_0_1_15_7: FA PORT MAP (CARRY_OUT_7(14),PARTIAL_PRODUCT_0_6(15),PARTIAL_PRODUCT_1_6(15),PARTIAL_PRODUCT_0_7(15),CARRY_OUT_7(15));
FA_C_0_1_16_7: FA PORT MAP (CARRY_OUT_7(15),PARTIAL_PRODUCT_0_6(16),PARTIAL_PRODUCT_1_6(16),PARTIAL_PRODUCT_0_7(16),CARRY_OUT_7(16));
FA_C_0_1_17_7: FA PORT MAP (CARRY_OUT_7(16),PARTIAL_PRODUCT_0_6(17),PARTIAL_PRODUCT_1_6(17),PARTIAL_PRODUCT_0_7(17),CARRY_OUT_7(17));
FA_C_0_1_18_7: FA PORT MAP (CARRY_OUT_7(17),PARTIAL_PRODUCT_0_6(18),PARTIAL_PRODUCT_1_6(18),PARTIAL_PRODUCT_0_7(18),CARRY_OUT_7(18));
FA_C_0_1_19_7: FA PORT MAP (CARRY_OUT_7(18),PARTIAL_PRODUCT_0_6(19),PARTIAL_PRODUCT_1_6(19),PARTIAL_PRODUCT_0_7(19),CARRY_OUT_7(19));
FA_C_0_1_20_7: FA PORT MAP (CARRY_OUT_7(19),PARTIAL_PRODUCT_0_6(20),PARTIAL_PRODUCT_1_6(20),PARTIAL_PRODUCT_0_7(20),CARRY_OUT_7(20));
FA_C_0_1_21_7: FA PORT MAP (CARRY_OUT_7(20),PARTIAL_PRODUCT_0_6(21),PARTIAL_PRODUCT_1_6(21),PARTIAL_PRODUCT_0_7(21),CARRY_OUT_7(21));
FA_C_0_1_22_7: FA PORT MAP (CARRY_OUT_7(21),PARTIAL_PRODUCT_0_6(22),PARTIAL_PRODUCT_1_6(22),PARTIAL_PRODUCT_0_7(22),CARRY_OUT_7(22));
FA_C_0_1_23_7: FA PORT MAP (CARRY_OUT_7(22),PARTIAL_PRODUCT_0_6(23),PARTIAL_PRODUCT_1_6(23),PARTIAL_PRODUCT_0_7(23),CARRY_OUT_7(23));
FA_C_0_1_24_7: FA PORT MAP (CARRY_OUT_7(23),PARTIAL_PRODUCT_0_6(24),PARTIAL_PRODUCT_1_6(24),PARTIAL_PRODUCT_0_7(24),CARRY_OUT_7(24));
FA_C_0_1_25_7: FA PORT MAP (CARRY_OUT_7(24),PARTIAL_PRODUCT_0_6(25),PARTIAL_PRODUCT_1_6(25),PARTIAL_PRODUCT_0_7(25),CARRY_OUT_7(25));
FA_C_0_1_26_7: FA PORT MAP (CARRY_OUT_7(25),PARTIAL_PRODUCT_0_6(26),PARTIAL_PRODUCT_1_6(26),PARTIAL_PRODUCT_0_7(26),CARRY_OUT_7(26));
FA_C_0_1_27_7: FA PORT MAP (CARRY_OUT_7(26),PARTIAL_PRODUCT_0_6(27),PARTIAL_PRODUCT_1_6(27),PARTIAL_PRODUCT_0_7(27),CARRY_OUT_7(27));
FA_C_0_1_28_7: FA PORT MAP (CARRY_OUT_7(27),PARTIAL_PRODUCT_0_6(28),PARTIAL_PRODUCT_1_6(28),PARTIAL_PRODUCT_0_7(28),CARRY_OUT_7(28));
FA_C_0_1_29_7: FA PORT MAP (CARRY_OUT_7(28),PARTIAL_PRODUCT_0_6(29),PARTIAL_PRODUCT_1_6(29),PARTIAL_PRODUCT_0_7(29),CARRY_OUT_7(29));
FA_C_0_1_30_7: FA PORT MAP (CARRY_OUT_7(29),PARTIAL_PRODUCT_0_6(30),PARTIAL_PRODUCT_1_6(30),PARTIAL_PRODUCT_0_7(30),CARRY_OUT_7(30));
FA_C_0_1_31_7: FA PORT MAP (CARRY_OUT_7(30),PARTIAL_PRODUCT_0_6(31),PARTIAL_PRODUCT_1_6(31),PARTIAL_PRODUCT_0_7(31),CARRY_OUT_7(31));
FA_C_0_1_32_7: FA PORT MAP (CARRY_OUT_7(31),PARTIAL_PRODUCT_0_6(32),PARTIAL_PRODUCT_1_6(32),PARTIAL_PRODUCT_0_7(32),CARRY_OUT_7(32));
FA_C_0_1_33_7: FA PORT MAP (CARRY_OUT_7(32),PARTIAL_PRODUCT_0_6(33),PARTIAL_PRODUCT_1_6(33),PARTIAL_PRODUCT_0_7(33),CARRY_OUT_7(33));
FA_C_0_1_34_7: FA PORT MAP (CARRY_OUT_7(33),PARTIAL_PRODUCT_0_6(34),PARTIAL_PRODUCT_1_6(34),PARTIAL_PRODUCT_0_7(34),CARRY_OUT_7(34));
FA_C_0_1_35_7: FA PORT MAP (CARRY_OUT_7(34),PARTIAL_PRODUCT_0_6(35),PARTIAL_PRODUCT_1_6(35),PARTIAL_PRODUCT_0_7(35),CARRY_OUT_7(35));
FA_C_0_1_36_7: FA PORT MAP (CARRY_OUT_7(35),PARTIAL_PRODUCT_0_6(36),PARTIAL_PRODUCT_1_6(36),PARTIAL_PRODUCT_0_7(36),CARRY_OUT_7(36));
FA_C_0_1_37_7: FA PORT MAP (CARRY_OUT_7(36),PARTIAL_PRODUCT_0_6(37),PARTIAL_PRODUCT_1_6(37),PARTIAL_PRODUCT_0_7(37),CARRY_OUT_7(37));
FA_C_0_1_38_7: FA PORT MAP (CARRY_OUT_7(37),PARTIAL_PRODUCT_0_6(38),PARTIAL_PRODUCT_1_6(38),PARTIAL_PRODUCT_0_7(38),CARRY_OUT_7(38));
FA_C_0_1_39_7: FA PORT MAP (CARRY_OUT_7(38),PARTIAL_PRODUCT_0_6(39),PARTIAL_PRODUCT_1_6(39),PARTIAL_PRODUCT_0_7(39),CARRY_OUT_7(39));
FA_C_0_1_40_7: FA PORT MAP (CARRY_OUT_7(39),PARTIAL_PRODUCT_0_6(40),PARTIAL_PRODUCT_1_6(40),PARTIAL_PRODUCT_0_7(40),CARRY_OUT_7(40));
FA_C_0_1_41_7: FA PORT MAP (CARRY_OUT_7(40),PARTIAL_PRODUCT_0_6(41),PARTIAL_PRODUCT_1_6(41),PARTIAL_PRODUCT_0_7(41),CARRY_OUT_7(41));
FA_C_0_1_42_7: FA PORT MAP (CARRY_OUT_7(41),PARTIAL_PRODUCT_0_6(42),PARTIAL_PRODUCT_1_6(42),PARTIAL_PRODUCT_0_7(42),CARRY_OUT_7(42));
FA_C_0_1_43_7: FA PORT MAP (CARRY_OUT_7(42),PARTIAL_PRODUCT_0_6(43),PARTIAL_PRODUCT_1_6(43),PARTIAL_PRODUCT_0_7(43),CARRY_OUT_7(43));
FA_C_0_1_44_7: FA PORT MAP (CARRY_OUT_7(43),PARTIAL_PRODUCT_0_6(44),PARTIAL_PRODUCT_1_6(44),PARTIAL_PRODUCT_0_7(44),CARRY_OUT_7(44));
FA_C_0_1_45_7: FA PORT MAP (CARRY_OUT_7(44),PARTIAL_PRODUCT_0_6(45),PARTIAL_PRODUCT_1_6(45),PARTIAL_PRODUCT_0_7(45),CARRY_OUT_7(45));
FA_C_0_1_46_7: FA PORT MAP (CARRY_OUT_7(45),PARTIAL_PRODUCT_0_6(46),PARTIAL_PRODUCT_1_6(46),PARTIAL_PRODUCT_0_7(46),CARRY_OUT_7(46));
FA_C_0_1_47_7: FA PORT MAP (CARRY_OUT_7(46),PARTIAL_PRODUCT_0_6(47),PARTIAL_PRODUCT_1_6(47),PARTIAL_PRODUCT_0_7(47),CARRY_OUT_7(47));
FA_C_0_1_48_7: FA PORT MAP (CARRY_OUT_7(47),PARTIAL_PRODUCT_0_6(48),PARTIAL_PRODUCT_1_6(48),PARTIAL_PRODUCT_0_7(48),CARRY_OUT_7(48));
FA_C_0_1_49_7: FA PORT MAP (CARRY_OUT_7(48),PARTIAL_PRODUCT_0_6(49),PARTIAL_PRODUCT_1_6(49),PARTIAL_PRODUCT_0_7(49),CARRY_OUT_7(49));
FA_C_0_1_50_7: FA PORT MAP (CARRY_OUT_7(49),PARTIAL_PRODUCT_0_6(50),PARTIAL_PRODUCT_1_6(50),PARTIAL_PRODUCT_0_7(50),CARRY_OUT_7(50));
FA_C_0_1_51_7: FA PORT MAP (CARRY_OUT_7(50),PARTIAL_PRODUCT_0_6(51),PARTIAL_PRODUCT_1_6(51),PARTIAL_PRODUCT_0_7(51),CARRY_OUT_7(51));
FA_C_0_1_52_7: FA PORT MAP (CARRY_OUT_7(51),PARTIAL_PRODUCT_0_6(52),PARTIAL_PRODUCT_1_6(52),PARTIAL_PRODUCT_0_7(52),CARRY_OUT_7(52));
FA_C_0_1_53_7: FA PORT MAP (CARRY_OUT_7(52),PARTIAL_PRODUCT_0_6(53),PARTIAL_PRODUCT_1_6(53),PARTIAL_PRODUCT_0_7(53),CARRY_OUT_7(53));
FA_C_0_1_54_7: FA PORT MAP (CARRY_OUT_7(53),PARTIAL_PRODUCT_0_6(54),PARTIAL_PRODUCT_1_6(54),PARTIAL_PRODUCT_0_7(54),CARRY_OUT_7(54));
FA_C_0_1_55_7: FA PORT MAP (CARRY_OUT_7(54),PARTIAL_PRODUCT_0_6(55),PARTIAL_PRODUCT_1_6(55),PARTIAL_PRODUCT_0_7(55),CARRY_OUT_7(55));
FA_C_0_1_56_7: FA PORT MAP (CARRY_OUT_7(55),PARTIAL_PRODUCT_0_6(56),PARTIAL_PRODUCT_1_6(56),PARTIAL_PRODUCT_0_7(56),CARRY_OUT_7(56));
FA_C_0_1_57_7: FA PORT MAP (CARRY_OUT_7(56),PARTIAL_PRODUCT_0_6(57),PARTIAL_PRODUCT_1_6(57),PARTIAL_PRODUCT_0_7(57),CARRY_OUT_7(57));
FA_C_0_1_58_7: FA PORT MAP (CARRY_OUT_7(57),PARTIAL_PRODUCT_0_6(58),PARTIAL_PRODUCT_1_6(58),PARTIAL_PRODUCT_0_7(58),CARRY_OUT_7(58));
FA_C_0_1_59_7: FA PORT MAP (CARRY_OUT_7(58),PARTIAL_PRODUCT_0_6(59),PARTIAL_PRODUCT_1_6(59),PARTIAL_PRODUCT_0_7(59),CARRY_OUT_7(59));
FA_C_0_1_60_7: FA PORT MAP (CARRY_OUT_7(59),PARTIAL_PRODUCT_0_6(60),PARTIAL_PRODUCT_1_6(60),PARTIAL_PRODUCT_0_7(60),CARRY_OUT_7(60));
FA_C_0_1_61_7: FA PORT MAP (CARRY_OUT_7(60),PARTIAL_PRODUCT_0_6(61),PARTIAL_PRODUCT_1_6(61),PARTIAL_PRODUCT_0_7(61),CARRY_OUT_7(61));
FA_C_0_1_62_7: FA PORT MAP (CARRY_OUT_7(61),PARTIAL_PRODUCT_0_6(62),PARTIAL_PRODUCT_1_6(62),PARTIAL_PRODUCT_0_7(62),CARRY_OUT_7(62));
FA_C_0_1_63_7: FA PORT MAP (CARRY_OUT_7(62),PARTIAL_PRODUCT_0_6(63),PARTIAL_PRODUCT_1_6(63),PARTIAL_PRODUCT_0_7(63),CARRY_OUT_7(63));


OUT_MULT <= PARTIAL_PRODUCT_0_7;


--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 6

--LEVEL 5 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 5

--LEVEL 4 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 4

--LEVEL 3 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 3

--LEVEL 2 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 2

--LEVEL 1 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 1

--LEVEL 0 DADDA TREE (COVER HA AND FA) --> HA_pp(i)_pp(i+1)_weight OR FA_pp(i)_pp(i+1)_pp(i+2)_weight <--

--NEW STRUCTURE OF PARTIAL PRODUCT PRODUCED BY LEVEL 0 --> FINAL RESULT

END ARCHITECTURE;


